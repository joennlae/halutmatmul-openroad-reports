module fp_16_32_adder__6142509188972423790 (operand_fp16_i,
    operand_fp32_i,
    result_o);
 input [15:0] operand_fp16_i;
 input [31:0] operand_fp32_i;
 output [31:0] result_o;

 wire _0000_;
 wire _0001_;
 wire net76;
 wire net75;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire net74;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire net73;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire net72;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire net71;
 wire _0024_;
 wire net70;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire net69;
 wire _0035_;
 wire net68;
 wire net67;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire net66;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire net65;
 wire net64;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire net63;
 wire _0067_;
 wire _0068_;
 wire net61;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire net60;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire net58;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire net57;
 wire net56;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire net54;
 wire net53;
 wire net52;
 wire _0130_;
 wire net51;
 wire net50;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire net49;
 wire _0139_;
 wire _0140_;
 wire net48;
 wire net47;
 wire net46;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire net45;
 wire net44;
 wire _0151_;
 wire net43;
 wire _0153_;
 wire _0154_;
 wire net42;
 wire net41;
 wire net40;
 wire _0158_;
 wire net39;
 wire net38;
 wire _0161_;
 wire net37;
 wire _0163_;
 wire _0164_;
 wire net36;
 wire net35;
 wire net34;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire net33;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire net32;
 wire net31;
 wire net30;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire net29;
 wire net28;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire net27;
 wire net26;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire net25;
 wire net24;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire net23;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire net22;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire net21;
 wire net20;
 wire _0276_;
 wire net19;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire net18;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire net17;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire net16;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire net15;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire net14;
 wire _0357_;
 wire net13;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire net11;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire net10;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire net9;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire net8;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire net7;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire net6;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire net5;
 wire net4;
 wire net3;
 wire net2;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire net1;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1079_;
 wire _1084_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1111_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1134_;
 wire _1135_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1196_;
 wire _1201_;
 wire _1202_;
 wire _1205_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1222_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1364_;
 wire _1365_;
 wire _1369_;
 wire net98;
 wire net97;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire net96;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire net95;
 wire _1388_;
 wire _1389_;
 wire net94;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire net93;
 wire net92;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire net91;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire net90;
 wire net89;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire net88;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire net87;
 wire _1439_;
 wire _1440_;
 wire net86;
 wire _1442_;
 wire net85;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire net84;
 wire _1456_;
 wire _1457_;
 wire net83;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire net82;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire net81;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire net80;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire net79;
 wire net78;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire net77;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire net62;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire net12;
 wire _1686_;
 wire _1687_;
 wire net55;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire net59;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1940_;
 wire _1941_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;

 BUF_X1 input41 (.A(operand_fp32_i[31]),
    .Z(net41));
 NOR2_X2 _1951_ (.A1(net4),
    .A2(net6),
    .ZN(_1071_));
 NOR3_X2 _1952_ (.A1(net3),
    .A2(net2),
    .A3(net5),
    .ZN(_1072_));
 AND2_X4 _1953_ (.A1(_1071_),
    .A2(_1072_),
    .ZN(_1073_));
 BUF_X1 input40 (.A(operand_fp32_i[30]),
    .Z(net40));
 BUF_X2 input39 (.A(operand_fp32_i[2]),
    .Z(net39));
 BUF_X2 input38 (.A(operand_fp32_i[29]),
    .Z(net38));
 BUF_X1 input37 (.A(operand_fp32_i[28]),
    .Z(net37));
 CLKBUF_X2 input36 (.A(operand_fp32_i[27]),
    .Z(net36));
 OR4_X4 _1959_ (.A1(net16),
    .A2(net15),
    .A3(net14),
    .A4(net13),
    .ZN(_1079_));
 BUF_X1 input35 (.A(operand_fp32_i[26]),
    .Z(net35));
 BUF_X2 input34 (.A(operand_fp32_i[25]),
    .Z(net34));
 BUF_X1 input33 (.A(operand_fp32_i[24]),
    .Z(net33));
 CLKBUF_X2 input32 (.A(operand_fp32_i[23]),
    .Z(net32));
 OR4_X2 _1964_ (.A1(net12),
    .A2(net11),
    .A3(net10),
    .A4(net9),
    .ZN(_1084_));
 BUF_X1 input31 (.A(operand_fp32_i[22]),
    .Z(net31));
 OR2_X2 _1966_ (.A1(net8),
    .A2(net1),
    .ZN(_1086_));
 NOR3_X2 _1967_ (.A1(_1079_),
    .A2(_1084_),
    .A3(_1086_),
    .ZN(_1087_));
 AOI21_X4 _1968_ (.A(net6),
    .B1(_1073_),
    .B2(_1087_),
    .ZN(_1540_));
 INV_X2 _1969_ (.A(_1540_),
    .ZN(_1535_));
 INV_X1 _1970_ (.A(net16),
    .ZN(_1088_));
 INV_X1 _1971_ (.A(net14),
    .ZN(_1089_));
 OAI21_X4 _1972_ (.A(_1088_),
    .B1(net15),
    .B2(_1089_),
    .ZN(_1090_));
 INV_X1 _1973_ (.A(net11),
    .ZN(_1091_));
 INV_X1 _1974_ (.A(net8),
    .ZN(_1092_));
 AOI21_X1 _1975_ (.A(net9),
    .B1(net1),
    .B2(_1092_),
    .ZN(_1093_));
 OAI21_X2 _1976_ (.A(_1091_),
    .B1(net10),
    .B2(_1093_),
    .ZN(_1094_));
 INV_X1 _1977_ (.A(net12),
    .ZN(_1095_));
 AOI21_X4 _1978_ (.A(_1079_),
    .B1(_1094_),
    .B2(_1095_),
    .ZN(_1096_));
 NOR2_X2 _1979_ (.A1(_1090_),
    .A2(_1096_),
    .ZN(_1799_));
 INV_X1 _1980_ (.A(_1799_),
    .ZN(_1803_));
 NOR4_X1 _1981_ (.A1(net12),
    .A2(net11),
    .A3(net10),
    .A4(net9),
    .ZN(_1097_));
 NOR3_X1 _1982_ (.A1(net12),
    .A2(net11),
    .A3(_1097_),
    .ZN(_1098_));
 NOR3_X1 _1983_ (.A1(net14),
    .A2(net13),
    .A3(_1098_),
    .ZN(_1099_));
 OR3_X1 _1984_ (.A1(net16),
    .A2(net15),
    .A3(_1099_),
    .ZN(_1804_));
 INV_X1 _1985_ (.A(_1804_),
    .ZN(_1800_));
 NAND2_X1 _1986_ (.A1(_1791_),
    .A2(_1079_),
    .ZN(_1100_));
 AOI21_X2 _1987_ (.A(net6),
    .B1(_1073_),
    .B2(_1100_),
    .ZN(_1527_));
 INV_X1 _1988_ (.A(_1527_),
    .ZN(_1531_));
 NOR4_X2 _1989_ (.A1(net16),
    .A2(net15),
    .A3(net14),
    .A4(net13),
    .ZN(_1101_));
 NAND2_X1 _1990_ (.A1(_1101_),
    .A2(_1084_),
    .ZN(_1792_));
 INV_X1 _1991_ (.A(_1792_),
    .ZN(_1810_));
 INV_X1 _1992_ (.A(net5),
    .ZN(_1102_));
 NAND2_X4 _1993_ (.A1(_1071_),
    .A2(_1072_),
    .ZN(_1103_));
 BUF_X1 input30 (.A(operand_fp32_i[21]),
    .Z(net30));
 NAND2_X1 _1995_ (.A1(_1793_),
    .A2(_1086_),
    .ZN(_1105_));
 NOR2_X1 _1996_ (.A1(_1079_),
    .A2(_1084_),
    .ZN(_1106_));
 MUX2_X1 _1997_ (.A(_1793_),
    .B(_1105_),
    .S(_1106_),
    .Z(_1107_));
 OAI21_X2 _1998_ (.A(_1102_),
    .B1(_1103_),
    .B2(_1107_),
    .ZN(_1785_));
 INV_X1 _1999_ (.A(_1785_),
    .ZN(_1788_));
 NOR2_X2 _2000_ (.A1(_1103_),
    .A2(_1087_),
    .ZN(_1108_));
 AOI21_X4 _2001_ (.A(net4),
    .B1(_1794_),
    .B2(_1108_),
    .ZN(_1519_));
 BUF_X1 input29 (.A(operand_fp32_i[20]),
    .Z(net29));
 BUF_X2 input28 (.A(operand_fp32_i[1]),
    .Z(net28));
 AOI21_X2 _2004_ (.A(net3),
    .B1(_1802_),
    .B2(_1108_),
    .ZN(_1511_));
 AOI21_X4 _2005_ (.A(net2),
    .B1(_1073_),
    .B2(_1799_),
    .ZN(_1843_));
 INV_X1 _2006_ (.A(net6),
    .ZN(_1768_));
 OR3_X1 _2007_ (.A1(_1079_),
    .A2(_1084_),
    .A3(_1086_),
    .ZN(_1111_));
 NOR2_X2 _2008_ (.A1(_1103_),
    .A2(_1111_),
    .ZN(_1807_));
 BUF_X1 input27 (.A(operand_fp32_i[19]),
    .Z(net27));
 AOI21_X1 _2010_ (.A(_1769_),
    .B1(_1773_),
    .B2(_1770_),
    .ZN(_1113_));
 OR2_X1 _2011_ (.A1(_1789_),
    .A2(_1797_),
    .ZN(_1114_));
 INV_X1 _2012_ (.A(_1517_),
    .ZN(_1115_));
 AOI21_X1 _2013_ (.A(_1114_),
    .B1(_1796_),
    .B2(_1115_),
    .ZN(_1116_));
 BUF_X1 input26 (.A(operand_fp32_i[18]),
    .Z(net26));
 AND4_X1 _2015_ (.A1(_1770_),
    .A2(_1777_),
    .A3(_1772_),
    .A4(_1781_),
    .ZN(_1118_));
 OR2_X1 _2016_ (.A1(_1787_),
    .A2(_1789_),
    .ZN(_1119_));
 NAND2_X1 _2017_ (.A1(_1118_),
    .A2(_1119_),
    .ZN(_1120_));
 NAND2_X1 _2018_ (.A1(_1770_),
    .A2(_1772_),
    .ZN(_1121_));
 AOI21_X1 _2019_ (.A(_1778_),
    .B1(_1782_),
    .B2(_1777_),
    .ZN(_1122_));
 OAI221_X2 _2020_ (.A(_1113_),
    .B1(_1116_),
    .B2(_1120_),
    .C1(_1121_),
    .C2(_1122_),
    .ZN(_1123_));
 BUF_X1 input25 (.A(operand_fp32_i[17]),
    .Z(net25));
 AND2_X1 _2022_ (.A1(_1518_),
    .A2(net92),
    .ZN(_1125_));
 OAI21_X1 _2023_ (.A(_1113_),
    .B1(_1121_),
    .B2(_1122_),
    .ZN(_1126_));
 NOR2_X1 _2024_ (.A1(_1789_),
    .A2(_1797_),
    .ZN(_1127_));
 INV_X1 _2025_ (.A(_1796_),
    .ZN(_1128_));
 OAI21_X2 _2026_ (.A(_1127_),
    .B1(_1128_),
    .B2(_1517_),
    .ZN(_1129_));
 AND2_X1 _2027_ (.A1(_1118_),
    .A2(_1119_),
    .ZN(_1130_));
 AOI21_X4 _2028_ (.A(_1126_),
    .B1(_1129_),
    .B2(_1130_),
    .ZN(_1131_));
 BUF_X1 input24 (.A(operand_fp32_i[16]),
    .Z(net24));
 BUF_X1 input23 (.A(operand_fp32_i[15]),
    .Z(net23));
 AOI21_X4 _2031_ (.A(_1125_),
    .B1(_1131_),
    .B2(_1513_),
    .ZN(_1134_));
 INV_X8 _2032_ (.A(_1134_),
    .ZN(_1135_));
 BUF_X1 input22 (.A(operand_fp32_i[14]),
    .Z(net22));
 BUF_X1 input21 (.A(operand_fp32_i[13]),
    .Z(net21));
 AND2_X1 _2035_ (.A1(_1525_),
    .A2(_1123_),
    .ZN(_1137_));
 AOI21_X4 _2036_ (.A(_1137_),
    .B1(_1131_),
    .B2(_1521_),
    .ZN(_1138_));
 INV_X8 _2037_ (.A(_1138_),
    .ZN(_1139_));
 CLKBUF_X2 input20 (.A(operand_fp32_i[12]),
    .Z(net20));
 CLKBUF_X2 input19 (.A(operand_fp32_i[11]),
    .Z(net19));
 BUF_X2 input18 (.A(operand_fp32_i[10]),
    .Z(net18));
 MUX2_X2 _2041_ (.A(_1530_),
    .B(_1534_),
    .S(_1123_),
    .Z(_1142_));
 INV_X2 _2042_ (.A(_1142_),
    .ZN(_1947_));
 INV_X1 _2043_ (.A(_1786_),
    .ZN(_1143_));
 INV_X1 _2044_ (.A(_1512_),
    .ZN(_1144_));
 AOI21_X1 _2045_ (.A(_1795_),
    .B1(_1796_),
    .B2(_1144_),
    .ZN(_1145_));
 INV_X1 _2046_ (.A(_1787_),
    .ZN(_1146_));
 OAI21_X1 _2047_ (.A(_1143_),
    .B1(_1145_),
    .B2(_1146_),
    .ZN(_1528_));
 AOI21_X1 _2048_ (.A(_1780_),
    .B1(_1528_),
    .B2(_1781_),
    .ZN(_1147_));
 INV_X1 _2049_ (.A(_1147_),
    .ZN(_1148_));
 AOI21_X1 _2050_ (.A(_1776_),
    .B1(_1148_),
    .B2(_1777_),
    .ZN(_1536_));
 INV_X1 _2051_ (.A(_1789_),
    .ZN(_1149_));
 AOI21_X1 _2052_ (.A(_1797_),
    .B1(_1796_),
    .B2(_1115_),
    .ZN(_1150_));
 OAI21_X1 _2053_ (.A(_1149_),
    .B1(_1150_),
    .B2(_1146_),
    .ZN(_1532_));
 AOI21_X1 _2054_ (.A(_1782_),
    .B1(_1532_),
    .B2(_1781_),
    .ZN(_1151_));
 INV_X1 _2055_ (.A(_1151_),
    .ZN(_1152_));
 AOI21_X1 _2056_ (.A(_1778_),
    .B1(_1152_),
    .B2(_1777_),
    .ZN(_1541_));
 MUX2_X2 _2057_ (.A(_1543_),
    .B(_1538_),
    .S(_1131_),
    .Z(_1930_));
 BUF_X2 input17 (.A(operand_fp32_i[0]),
    .Z(net17));
 NAND3_X1 _2059_ (.A1(_1815_),
    .A2(_1809_),
    .A3(_1818_),
    .ZN(_1154_));
 INV_X1 _2060_ (.A(_1823_),
    .ZN(_1155_));
 AOI21_X1 _2061_ (.A(_1826_),
    .B1(_1827_),
    .B2(_1829_),
    .ZN(_1156_));
 INV_X1 _2062_ (.A(_1824_),
    .ZN(_1157_));
 OAI21_X1 _2063_ (.A(_1155_),
    .B1(_1156_),
    .B2(_1157_),
    .ZN(_1158_));
 AOI21_X1 _2064_ (.A(_1820_),
    .B1(_1158_),
    .B2(_1821_),
    .ZN(_1159_));
 NAND4_X1 _2065_ (.A1(_1821_),
    .A2(_1824_),
    .A3(_1827_),
    .A4(_1830_),
    .ZN(_1160_));
 AOI21_X1 _2066_ (.A(_1154_),
    .B1(_1159_),
    .B2(_1160_),
    .ZN(_1161_));
 AND2_X1 _2067_ (.A1(_1833_),
    .A2(_1161_),
    .ZN(_1162_));
 INV_X1 _2068_ (.A(_1836_),
    .ZN(_1163_));
 INV_X1 _2069_ (.A(_1838_),
    .ZN(_1164_));
 BUF_X4 input16 (.A(operand_fp16_i[9]),
    .Z(net16));
 NAND4_X1 _2071_ (.A1(_1811_),
    .A2(_1101_),
    .A3(_1097_),
    .A4(_1086_),
    .ZN(_1166_));
 OAI21_X1 _2072_ (.A(_1166_),
    .B1(_1106_),
    .B2(_1811_),
    .ZN(_1167_));
 NAND2_X1 _2073_ (.A1(_1073_),
    .A2(_1167_),
    .ZN(_1168_));
 NOR2_X1 _2074_ (.A1(_1812_),
    .A2(_1168_),
    .ZN(_1169_));
 INV_X1 _2075_ (.A(net1),
    .ZN(_1170_));
 NOR4_X4 _2076_ (.A1(_1170_),
    .A2(net98),
    .A3(_1090_),
    .A4(_1096_),
    .ZN(_1171_));
 AOI22_X4 _2077_ (.A1(net1),
    .A2(_1103_),
    .B1(_1169_),
    .B2(_1171_),
    .ZN(_1172_));
 OAI21_X1 _2078_ (.A(_1839_),
    .B1(_1172_),
    .B2(net21),
    .ZN(_1173_));
 AOI21_X1 _2079_ (.A(_1163_),
    .B1(_1164_),
    .B2(_1173_),
    .ZN(_1174_));
 OAI21_X2 _2080_ (.A(_1162_),
    .B1(_1174_),
    .B2(_1835_),
    .ZN(_1175_));
 INV_X1 _2081_ (.A(_1808_),
    .ZN(_1176_));
 AND2_X1 _2082_ (.A1(_1815_),
    .A2(_1817_),
    .ZN(_1177_));
 OAI21_X1 _2083_ (.A(_1809_),
    .B1(_1814_),
    .B2(_1177_),
    .ZN(_1178_));
 INV_X1 _2084_ (.A(_1159_),
    .ZN(_1179_));
 OAI21_X1 _2085_ (.A(_1161_),
    .B1(_1179_),
    .B2(_1832_),
    .ZN(_1180_));
 AND4_X1 _2086_ (.A1(_1176_),
    .A2(_1940_),
    .A3(_1178_),
    .A4(_1180_),
    .ZN(_1181_));
 MUX2_X2 _2087_ (.A(_1537_),
    .B(_1542_),
    .S(_1123_),
    .Z(_1182_));
 XOR2_X2 _2088_ (.A(_1770_),
    .B(_1182_),
    .Z(_1183_));
 AND2_X4 _2089_ (.A1(_1930_),
    .A2(_1183_),
    .ZN(_1184_));
 NAND2_X2 _2090_ (.A1(_1139_),
    .A2(_1184_),
    .ZN(_1185_));
 MUX2_X2 _2091_ (.A(_1520_),
    .B(_1524_),
    .S(_1123_),
    .Z(_1186_));
 XNOR2_X2 _2092_ (.A(_1146_),
    .B(_1186_),
    .ZN(_1187_));
 MUX2_X2 _2093_ (.A(_1529_),
    .B(_1533_),
    .S(net92),
    .Z(_1188_));
 XOR2_X2 _2094_ (.A(_1777_),
    .B(_1188_),
    .Z(_1189_));
 NOR2_X4 _2095_ (.A1(_1947_),
    .A2(_1189_),
    .ZN(_1190_));
 NAND2_X4 _2096_ (.A1(_1187_),
    .A2(_1190_),
    .ZN(_1191_));
 NOR2_X1 _2097_ (.A1(_1185_),
    .A2(_1191_),
    .ZN(_1192_));
 AND3_X1 _2098_ (.A1(_1175_),
    .A2(_1181_),
    .A3(_1192_),
    .ZN(_1193_));
 NOR2_X1 _2099_ (.A1(_1131_),
    .A2(_1193_),
    .ZN(_1194_));
 MUX2_X1 _2100_ (.A(net7),
    .B(net41),
    .S(_1194_),
    .Z(net73));
 CLKBUF_X3 input15 (.A(operand_fp16_i[8]),
    .Z(net15));
 INV_X8 _2102_ (.A(net95),
    .ZN(_1196_));
 BUF_X4 input14 (.A(operand_fp16_i[7]),
    .Z(net14));
 CLKBUF_X3 input13 (.A(operand_fp16_i[6]),
    .Z(net13));
 CLKBUF_X3 input12 (.A(operand_fp16_i[5]),
    .Z(net12));
 BUF_X2 input11 (.A(operand_fp16_i[4]),
    .Z(net11));
 XOR2_X2 _2107_ (.A(net7),
    .B(net41),
    .Z(_1613_));
 CLKBUF_X2 input10 (.A(operand_fp16_i[3]),
    .Z(net10));
 BUF_X1 input9 (.A(operand_fp16_i[2]),
    .Z(net9));
 NAND4_X4 _2110_ (.A1(net91),
    .A2(_1175_),
    .A3(_1181_),
    .A4(_1192_),
    .ZN(_1201_));
 NAND2_X4 _2111_ (.A1(_1613_),
    .A2(_1201_),
    .ZN(_1202_));
 BUF_X1 input8 (.A(operand_fp16_i[1]),
    .Z(net8));
 BUF_X1 input7 (.A(operand_fp16_i[15]),
    .Z(net7));
 XNOR2_X2 _2114_ (.A(_1787_),
    .B(_1186_),
    .ZN(_1205_));
 CLKBUF_X3 input6 (.A(operand_fp16_i[14]),
    .Z(net6));
 XNOR2_X2 _2116_ (.A(_1777_),
    .B(_1188_),
    .ZN(_1207_));
 NAND2_X2 _2117_ (.A1(_1142_),
    .A2(_1207_),
    .ZN(_1208_));
 NOR2_X4 _2118_ (.A1(_1205_),
    .A2(_1208_),
    .ZN(_1209_));
 BUF_X1 input5 (.A(operand_fp16_i[13]),
    .Z(net5));
 CLKBUF_X2 input4 (.A(operand_fp16_i[12]),
    .Z(net4));
 BUF_X1 input3 (.A(operand_fp16_i[11]),
    .Z(net3));
 CLKBUF_X2 input2 (.A(operand_fp16_i[10]),
    .Z(net2));
 NOR4_X1 _2123_ (.A1(net37),
    .A2(net36),
    .A3(net40),
    .A4(net38),
    .ZN(_1214_));
 NOR4_X1 _2124_ (.A1(net33),
    .A2(net32),
    .A3(net35),
    .A4(net34),
    .ZN(_1215_));
 NAND2_X1 _2125_ (.A1(_1214_),
    .A2(_1215_),
    .ZN(_1806_));
 NOR2_X1 _2126_ (.A1(net92),
    .A2(_1806_),
    .ZN(_1216_));
 AOI21_X2 _2127_ (.A(_1216_),
    .B1(net92),
    .B2(_1807_),
    .ZN(_1217_));
 NAND2_X1 _2128_ (.A1(_1842_),
    .A2(_1217_),
    .ZN(_1218_));
 NOR3_X2 _2129_ (.A1(_1134_),
    .A2(_1185_),
    .A3(_1218_),
    .ZN(_1219_));
 NAND2_X1 _2130_ (.A1(_1209_),
    .A2(_1219_),
    .ZN(_1220_));
 XNOR2_X1 _2131_ (.A(_1202_),
    .B(_1220_),
    .ZN(_1546_));
 CLKBUF_X3 input1 (.A(operand_fp16_i[0]),
    .Z(net1));
 AND3_X4 _2133_ (.A1(net92),
    .A2(_1193_),
    .A3(_1613_),
    .ZN(_1222_));
 TAPCELL_X1 PHY_109 ();
 TAPCELL_X1 PHY_108 ();
 TAPCELL_X1 PHY_107 ();
 NAND2_X1 _2137_ (.A1(_1807_),
    .A2(_1131_),
    .ZN(_1225_));
 OAI21_X1 _2138_ (.A(_1225_),
    .B1(_1806_),
    .B2(_1131_),
    .ZN(_1226_));
 XOR2_X2 _2139_ (.A(_1222_),
    .B(_1226_),
    .Z(_1545_));
 INV_X1 _2140_ (.A(_1812_),
    .ZN(_1227_));
 NAND2_X1 _2141_ (.A1(_1106_),
    .A2(_1086_),
    .ZN(_1228_));
 XOR2_X2 _2142_ (.A(_1811_),
    .B(_1228_),
    .Z(_1229_));
 OAI21_X2 _2143_ (.A(net1),
    .B1(_1090_),
    .B2(_1096_),
    .ZN(_1230_));
 INV_X1 _2144_ (.A(net15),
    .ZN(_1231_));
 AOI21_X4 _2145_ (.A(net16),
    .B1(_1231_),
    .B2(net14),
    .ZN(_1232_));
 INV_X1 _2146_ (.A(net10),
    .ZN(_1233_));
 INV_X1 _2147_ (.A(net9),
    .ZN(_1234_));
 OAI21_X1 _2148_ (.A(_1234_),
    .B1(_1170_),
    .B2(net8),
    .ZN(_1235_));
 AOI21_X1 _2149_ (.A(net11),
    .B1(_1233_),
    .B2(_1235_),
    .ZN(_1236_));
 OAI21_X2 _2150_ (.A(_1101_),
    .B1(_1236_),
    .B2(net12),
    .ZN(_1237_));
 NAND3_X2 _2151_ (.A1(net8),
    .A2(_1232_),
    .A3(_1237_),
    .ZN(_1238_));
 AOI211_X2 _2152_ (.A(_1802_),
    .B(_1229_),
    .C1(_1230_),
    .C2(_1238_),
    .ZN(_1239_));
 INV_X1 _2153_ (.A(_1229_),
    .ZN(_1240_));
 INV_X2 _2154_ (.A(_1802_),
    .ZN(_1241_));
 AOI21_X1 _2155_ (.A(net13),
    .B1(net15),
    .B2(_1088_),
    .ZN(_1242_));
 NOR3_X1 _2156_ (.A1(_1089_),
    .A2(_1241_),
    .A3(_1242_),
    .ZN(_1243_));
 MUX2_X1 _2157_ (.A(net15),
    .B(net13),
    .S(_1802_),
    .Z(_1244_));
 AOI21_X1 _2158_ (.A(_1243_),
    .B1(_1244_),
    .B2(net16),
    .ZN(_1245_));
 NOR2_X1 _2159_ (.A1(_1240_),
    .A2(_1245_),
    .ZN(_1246_));
 OAI21_X1 _2160_ (.A(_1227_),
    .B1(_1239_),
    .B2(_1246_),
    .ZN(_1247_));
 NAND2_X1 _2161_ (.A1(_1812_),
    .A2(_1229_),
    .ZN(_1248_));
 INV_X1 _2162_ (.A(_1248_),
    .ZN(_1249_));
 NAND2_X1 _2163_ (.A1(_1079_),
    .A2(_1232_),
    .ZN(_1250_));
 AOI22_X1 _2164_ (.A1(_1095_),
    .A2(_1232_),
    .B1(_1250_),
    .B2(_1091_),
    .ZN(_1251_));
 INV_X1 _2165_ (.A(_1251_),
    .ZN(_1252_));
 NOR2_X1 _2166_ (.A1(_1802_),
    .A2(_1252_),
    .ZN(_1253_));
 NAND3_X1 _2167_ (.A1(net10),
    .A2(_1232_),
    .A3(_1237_),
    .ZN(_1254_));
 OAI21_X1 _2168_ (.A(net9),
    .B1(_1090_),
    .B2(_1096_),
    .ZN(_1255_));
 AOI21_X1 _2169_ (.A(_1241_),
    .B1(_1254_),
    .B2(_1255_),
    .ZN(_1256_));
 OAI21_X1 _2170_ (.A(_1249_),
    .B1(_1253_),
    .B2(_1256_),
    .ZN(_1257_));
 AOI21_X1 _2171_ (.A(_1103_),
    .B1(_1247_),
    .B2(_1257_),
    .ZN(_1258_));
 AOI21_X1 _2172_ (.A(_1258_),
    .B1(_1103_),
    .B2(net16),
    .ZN(_1813_));
 NOR2_X1 _2173_ (.A1(_1171_),
    .A2(_1229_),
    .ZN(_1259_));
 NAND3_X1 _2174_ (.A1(_1089_),
    .A2(net13),
    .A3(_1802_),
    .ZN(_1260_));
 OAI21_X1 _2175_ (.A(net15),
    .B1(net13),
    .B2(_1241_),
    .ZN(_1261_));
 AOI21_X1 _2176_ (.A(net16),
    .B1(_1260_),
    .B2(_1261_),
    .ZN(_1262_));
 AOI21_X1 _2177_ (.A(_1095_),
    .B1(net15),
    .B2(_1088_),
    .ZN(_1263_));
 MUX2_X1 _2178_ (.A(net14),
    .B(_1263_),
    .S(_1802_),
    .Z(_1264_));
 NOR3_X1 _2179_ (.A1(_1240_),
    .A2(_1262_),
    .A3(_1264_),
    .ZN(_1265_));
 NAND2_X1 _2180_ (.A1(net10),
    .A2(_1250_),
    .ZN(_1266_));
 NAND2_X1 _2181_ (.A1(net12),
    .A2(_1101_),
    .ZN(_1267_));
 NAND3_X1 _2182_ (.A1(net11),
    .A2(_1232_),
    .A3(_1267_),
    .ZN(_1268_));
 NAND2_X1 _2183_ (.A1(_1266_),
    .A2(_1268_),
    .ZN(_1269_));
 NOR2_X1 _2184_ (.A1(net98),
    .A2(_1269_),
    .ZN(_1270_));
 NOR3_X1 _2185_ (.A1(_1234_),
    .A2(_1090_),
    .A3(_1096_),
    .ZN(_1271_));
 AOI21_X1 _2186_ (.A(_1092_),
    .B1(_1232_),
    .B2(_1237_),
    .ZN(_1272_));
 NOR3_X1 _2187_ (.A1(_1241_),
    .A2(_1271_),
    .A3(_1272_),
    .ZN(_1273_));
 OAI33_X1 _2188_ (.A1(_1812_),
    .A2(_1259_),
    .A3(_1265_),
    .B1(_1270_),
    .B2(_1273_),
    .B3(_1248_),
    .ZN(_1274_));
 MUX2_X1 _2189_ (.A(net15),
    .B(_1274_),
    .S(_1073_),
    .Z(_1275_));
 INV_X1 _2190_ (.A(_1275_),
    .ZN(_1816_));
 AND2_X2 _2191_ (.A1(_1073_),
    .A2(_1167_),
    .ZN(_1276_));
 OAI21_X1 _2192_ (.A(_1241_),
    .B1(net14),
    .B2(net16),
    .ZN(_1277_));
 OAI22_X1 _2193_ (.A1(_1241_),
    .A2(_1252_),
    .B1(_1277_),
    .B2(_1242_),
    .ZN(_1278_));
 NOR2_X1 _2194_ (.A1(_1812_),
    .A2(_1278_),
    .ZN(_1279_));
 NAND3_X1 _2195_ (.A1(net98),
    .A2(_1238_),
    .A3(_1230_),
    .ZN(_1280_));
 NAND2_X1 _2196_ (.A1(_1254_),
    .A2(_1255_),
    .ZN(_1281_));
 OAI21_X2 _2197_ (.A(_1280_),
    .B1(_1281_),
    .B2(net98),
    .ZN(_1282_));
 AOI21_X2 _2198_ (.A(_1279_),
    .B1(_1282_),
    .B2(_1812_),
    .ZN(_1283_));
 AOI22_X4 _2199_ (.A1(net14),
    .A2(_1103_),
    .B1(_1276_),
    .B2(_1283_),
    .ZN(_1819_));
 AND2_X1 _2200_ (.A1(net13),
    .A2(_1103_),
    .ZN(_1284_));
 NOR3_X1 _2201_ (.A1(net98),
    .A2(_1271_),
    .A3(_1272_),
    .ZN(_1285_));
 AOI21_X1 _2202_ (.A(_1241_),
    .B1(_1799_),
    .B2(net1),
    .ZN(_1286_));
 OR2_X1 _2203_ (.A1(_1285_),
    .A2(_1286_),
    .ZN(_1287_));
 AOI22_X1 _2204_ (.A1(net13),
    .A2(_1232_),
    .B1(_1250_),
    .B2(net12),
    .ZN(_1288_));
 NOR2_X1 _2205_ (.A1(net98),
    .A2(_1288_),
    .ZN(_1289_));
 AOI21_X1 _2206_ (.A(_1289_),
    .B1(_1269_),
    .B2(net98),
    .ZN(_1290_));
 MUX2_X1 _2207_ (.A(_1287_),
    .B(_1290_),
    .S(_1227_),
    .Z(_1291_));
 NOR2_X1 _2208_ (.A1(_1168_),
    .A2(_1291_),
    .ZN(_1292_));
 NOR2_X1 _2209_ (.A1(_1284_),
    .A2(_1292_),
    .ZN(_1822_));
 NAND2_X1 _2210_ (.A1(_1238_),
    .A2(_1230_),
    .ZN(_1293_));
 NAND2_X1 _2211_ (.A1(_1241_),
    .A2(_1293_),
    .ZN(_1294_));
 NOR2_X1 _2212_ (.A1(_1256_),
    .A2(_1253_),
    .ZN(_1295_));
 MUX2_X1 _2213_ (.A(_1294_),
    .B(_1295_),
    .S(_1227_),
    .Z(_1296_));
 NOR2_X1 _2214_ (.A1(_1168_),
    .A2(_1296_),
    .ZN(_1297_));
 AOI21_X1 _2215_ (.A(_1297_),
    .B1(_1103_),
    .B2(net12),
    .ZN(_1825_));
 NAND2_X1 _2216_ (.A1(net11),
    .A2(_1103_),
    .ZN(_1298_));
 AND2_X1 _2217_ (.A1(_1812_),
    .A2(_1171_),
    .ZN(_1299_));
 NOR3_X1 _2218_ (.A1(_1812_),
    .A2(_1270_),
    .A3(_1273_),
    .ZN(_1300_));
 OAI21_X1 _2219_ (.A(_1276_),
    .B1(_1299_),
    .B2(_1300_),
    .ZN(_1301_));
 AND2_X1 _2220_ (.A1(_1298_),
    .A2(_1301_),
    .ZN(_1828_));
 NAND2_X2 _2221_ (.A1(_1227_),
    .A2(_1276_),
    .ZN(_1302_));
 OAI22_X4 _2222_ (.A1(_1233_),
    .A2(_1073_),
    .B1(_1302_),
    .B2(_1282_),
    .ZN(_1303_));
 INV_X1 _2223_ (.A(_1303_),
    .ZN(_1831_));
 OAI22_X1 _2224_ (.A1(_1234_),
    .A2(_1073_),
    .B1(_1302_),
    .B2(_1287_),
    .ZN(_1304_));
 INV_X1 _2225_ (.A(_1304_),
    .ZN(_1834_));
 AOI211_X2 _2226_ (.A(net98),
    .B(_1302_),
    .C1(_1238_),
    .C2(_1230_),
    .ZN(_1305_));
 NOR2_X1 _2227_ (.A1(_1092_),
    .A2(_1073_),
    .ZN(_1306_));
 NOR2_X1 _2228_ (.A1(_1305_),
    .A2(_1306_),
    .ZN(_1837_));
 NAND2_X4 _2229_ (.A1(_1205_),
    .A2(_1190_),
    .ZN(_1307_));
 AND2_X1 _2230_ (.A1(net30),
    .A2(_1131_),
    .ZN(_1308_));
 AOI21_X2 _2231_ (.A(_1308_),
    .B1(_1275_),
    .B2(net92),
    .ZN(_1309_));
 AOI21_X1 _2232_ (.A(_1131_),
    .B1(_1103_),
    .B2(net16),
    .ZN(_1310_));
 INV_X1 _2233_ (.A(net31),
    .ZN(_1311_));
 AOI21_X1 _2234_ (.A(_1310_),
    .B1(_1131_),
    .B2(_1311_),
    .ZN(_1312_));
 AOI21_X1 _2235_ (.A(_1312_),
    .B1(_1258_),
    .B2(net92),
    .ZN(_1313_));
 MUX2_X1 _2236_ (.A(_1309_),
    .B(_1313_),
    .S(_1196_),
    .Z(_1314_));
 MUX2_X2 _2237_ (.A(_1218_),
    .B(_1314_),
    .S(_1135_),
    .Z(_1315_));
 NOR3_X1 _2238_ (.A1(_1185_),
    .A2(_1307_),
    .A3(_1315_),
    .ZN(_1316_));
 OR2_X1 _2239_ (.A1(net27),
    .A2(net90),
    .ZN(_1317_));
 NOR3_X1 _2240_ (.A1(_1227_),
    .A2(_1131_),
    .A3(_1284_),
    .ZN(_1318_));
 OAI21_X1 _2241_ (.A(_1318_),
    .B1(_1286_),
    .B2(_1285_),
    .ZN(_1319_));
 NOR3_X1 _2242_ (.A1(_1131_),
    .A2(_1276_),
    .A3(_1284_),
    .ZN(_1320_));
 NOR3_X1 _2243_ (.A1(_1812_),
    .A2(_1131_),
    .A3(_1284_),
    .ZN(_1321_));
 AOI21_X1 _2244_ (.A(_1320_),
    .B1(_1321_),
    .B2(_1290_),
    .ZN(_1322_));
 NAND3_X1 _2245_ (.A1(_1317_),
    .A2(_1319_),
    .A3(_1322_),
    .ZN(_1323_));
 NOR2_X1 _2246_ (.A1(_1196_),
    .A2(_1323_),
    .ZN(_1324_));
 INV_X1 _2247_ (.A(_1324_),
    .ZN(_1325_));
 INV_X1 _2248_ (.A(net29),
    .ZN(_1326_));
 MUX2_X1 _2249_ (.A(_1326_),
    .B(_1819_),
    .S(net90),
    .Z(_1327_));
 OAI21_X2 _2250_ (.A(_1325_),
    .B1(_1327_),
    .B2(net96),
    .ZN(_1328_));
 NOR2_X1 _2251_ (.A1(net25),
    .A2(net90),
    .ZN(_1329_));
 AND2_X1 _2252_ (.A1(net90),
    .A2(_1298_),
    .ZN(_1330_));
 AOI21_X2 _2253_ (.A(_1329_),
    .B1(_1330_),
    .B2(_1301_),
    .ZN(_1331_));
 NAND3_X1 _2254_ (.A1(net12),
    .A2(_1103_),
    .A3(net90),
    .ZN(_1332_));
 NAND2_X1 _2255_ (.A1(net90),
    .A2(_1276_),
    .ZN(_1333_));
 INV_X1 _2256_ (.A(net26),
    .ZN(_1334_));
 OAI221_X2 _2257_ (.A(_1332_),
    .B1(_1333_),
    .B2(_1296_),
    .C1(_1334_),
    .C2(net90),
    .ZN(_1335_));
 MUX2_X1 _2258_ (.A(_1331_),
    .B(_1335_),
    .S(_1196_),
    .Z(_1336_));
 TAPCELL_X1 PHY_106 ();
 MUX2_X1 _2260_ (.A(_1328_),
    .B(_1336_),
    .S(_1135_),
    .Z(_1338_));
 NAND2_X1 _2261_ (.A1(net21),
    .A2(_1131_),
    .ZN(_1339_));
 OAI21_X2 _2262_ (.A(_1339_),
    .B1(_1172_),
    .B2(_1131_),
    .ZN(_1340_));
 NAND2_X1 _2263_ (.A1(net96),
    .A2(_1340_),
    .ZN(_1341_));
 OR3_X1 _2264_ (.A1(_1131_),
    .A2(_1305_),
    .A3(_1306_),
    .ZN(_1342_));
 OR2_X1 _2265_ (.A1(net22),
    .A2(net90),
    .ZN(_1343_));
 NAND3_X1 _2266_ (.A1(_1196_),
    .A2(_1342_),
    .A3(_1343_),
    .ZN(_1344_));
 NAND3_X1 _2267_ (.A1(_1135_),
    .A2(_1341_),
    .A3(_1344_),
    .ZN(_1345_));
 OR2_X1 _2268_ (.A1(net23),
    .A2(net90),
    .ZN(_1346_));
 OAI221_X2 _2269_ (.A(net90),
    .B1(_1302_),
    .B2(_1287_),
    .C1(_1073_),
    .C2(_1234_),
    .ZN(_1347_));
 NAND3_X1 _2270_ (.A1(net96),
    .A2(_1346_),
    .A3(_1347_),
    .ZN(_1348_));
 OR2_X1 _2271_ (.A1(net24),
    .A2(net90),
    .ZN(_1349_));
 OAI21_X4 _2272_ (.A(_1349_),
    .B1(_1303_),
    .B2(_1131_),
    .ZN(_1350_));
 OAI21_X1 _2273_ (.A(_1348_),
    .B1(_1350_),
    .B2(net97),
    .ZN(_1351_));
 OR2_X1 _2274_ (.A1(_1135_),
    .A2(_1351_),
    .ZN(_1352_));
 AND2_X1 _2275_ (.A1(_1345_),
    .A2(_1352_),
    .ZN(_1353_));
 MUX2_X1 _2276_ (.A(_1338_),
    .B(_1353_),
    .S(_1139_),
    .Z(_1354_));
 NAND2_X4 _2277_ (.A1(_1930_),
    .A2(_1183_),
    .ZN(_1355_));
 TAPCELL_X1 PHY_105 ();
 TAPCELL_X1 PHY_104 ();
 NOR2_X1 _2280_ (.A1(_1355_),
    .A2(_1191_),
    .ZN(_1358_));
 AOI21_X1 _2281_ (.A(_1316_),
    .B1(_1354_),
    .B2(_1358_),
    .ZN(_1359_));
 XNOR2_X1 _2282_ (.A(_1202_),
    .B(_1359_),
    .ZN(_1571_));
 NAND2_X1 _2283_ (.A1(net21),
    .A2(net90),
    .ZN(_1360_));
 OAI21_X2 _2284_ (.A(_1360_),
    .B1(_1172_),
    .B2(net90),
    .ZN(_1361_));
 XOR2_X2 _2285_ (.A(_1222_),
    .B(_1361_),
    .Z(_1873_));
 INV_X1 _2286_ (.A(_1873_),
    .ZN(_1570_));
 NAND2_X1 _2287_ (.A1(_1190_),
    .A2(_1202_),
    .ZN(_1362_));
 TAPCELL_X1 PHY_103 ();
 AND3_X1 _2289_ (.A1(_1138_),
    .A2(_1184_),
    .A3(_1345_),
    .ZN(_1364_));
 NOR2_X4 _2290_ (.A1(net91),
    .A2(_1355_),
    .ZN(_1365_));
 TAPCELL_X1 PHY_102 ();
 TAPCELL_X1 PHY_101 ();
 TAPCELL_X1 PHY_100 ();
 MUX2_X1 _2294_ (.A(net20),
    .B(net19),
    .S(net97),
    .Z(_1369_));
 TAPCELL_X1 PHY_99 ();
 TAPCELL_X1 PHY_98 ();
 MUX2_X1 _2297_ (.A(net18),
    .B(net48),
    .S(net97),
    .Z(_1372_));
 MUX2_X1 _2298_ (.A(_1369_),
    .B(_1372_),
    .S(_1135_),
    .Z(_1373_));
 NAND2_X1 _2299_ (.A1(_1365_),
    .A2(_1373_),
    .ZN(_1374_));
 INV_X1 _2300_ (.A(_1374_),
    .ZN(_1375_));
 AOI22_X2 _2301_ (.A1(_1352_),
    .A2(_1364_),
    .B1(_1375_),
    .B2(_1139_),
    .ZN(_1376_));
 MUX2_X1 _2302_ (.A(_1362_),
    .B(_1202_),
    .S(_1376_),
    .Z(_1377_));
 OAI22_X1 _2303_ (.A1(_1190_),
    .A2(_1202_),
    .B1(_1377_),
    .B2(_1205_),
    .ZN(_1378_));
 AND2_X4 _2304_ (.A1(_1613_),
    .A2(_1201_),
    .ZN(_1379_));
 TAPCELL_X1 PHY_97 ();
 INV_X1 _2306_ (.A(_1362_),
    .ZN(_1381_));
 OR2_X1 _2307_ (.A1(_1134_),
    .A2(_1336_),
    .ZN(_1382_));
 OAI21_X2 _2308_ (.A(_1382_),
    .B1(_1328_),
    .B2(_1135_),
    .ZN(_1383_));
 NAND2_X2 _2309_ (.A1(_1138_),
    .A2(_1184_),
    .ZN(_1384_));
 OAI22_X4 _2310_ (.A1(_1185_),
    .A2(_1383_),
    .B1(_1315_),
    .B2(_1384_),
    .ZN(_1385_));
 MUX2_X1 _2311_ (.A(_1379_),
    .B(_1381_),
    .S(_1385_),
    .Z(_1386_));
 AOI21_X1 _2312_ (.A(_1378_),
    .B1(_1386_),
    .B2(_1205_),
    .ZN(_1581_));
 TAPCELL_X1 PHY_96 ();
 NAND2_X1 _2314_ (.A1(net48),
    .A2(net91),
    .ZN(_1388_));
 XNOR2_X1 _2315_ (.A(_1222_),
    .B(_1388_),
    .ZN(_1887_));
 INV_X1 _2316_ (.A(_1887_),
    .ZN(_1580_));
 NAND2_X1 _2317_ (.A1(_1142_),
    .A2(_1202_),
    .ZN(_1389_));
 TAPCELL_X1 PHY_95 ();
 AOI21_X1 _2319_ (.A(_1135_),
    .B1(_1341_),
    .B2(_1344_),
    .ZN(_1391_));
 AND3_X1 _2320_ (.A1(_1513_),
    .A2(_1131_),
    .A3(_1369_),
    .ZN(_1392_));
 OAI21_X1 _2321_ (.A(_1184_),
    .B1(_1391_),
    .B2(_1392_),
    .ZN(_1393_));
 TAPCELL_X1 PHY_94 ();
 TAPCELL_X1 PHY_93 ();
 MUX2_X1 _2324_ (.A(net47),
    .B(net46),
    .S(net94),
    .Z(_1396_));
 MUX2_X1 _2325_ (.A(_1372_),
    .B(_1396_),
    .S(_1135_),
    .Z(_1397_));
 NAND2_X1 _2326_ (.A1(_1365_),
    .A2(_1397_),
    .ZN(_1398_));
 MUX2_X1 _2327_ (.A(_1393_),
    .B(_1398_),
    .S(_1139_),
    .Z(_1399_));
 NAND2_X1 _2328_ (.A1(_1187_),
    .A2(_1399_),
    .ZN(_1400_));
 NAND3_X1 _2329_ (.A1(_1190_),
    .A2(_1379_),
    .A3(_1400_),
    .ZN(_1401_));
 NOR2_X2 _2330_ (.A1(_1138_),
    .A2(_1355_),
    .ZN(_1402_));
 OAI211_X2 _2331_ (.A(_1135_),
    .B(_1348_),
    .C1(_1350_),
    .C2(net97),
    .ZN(_1403_));
 OAI211_X2 _2332_ (.A(_1402_),
    .B(_1403_),
    .C1(_1336_),
    .C2(_1135_),
    .ZN(_1404_));
 AND2_X1 _2333_ (.A1(_1205_),
    .A2(_1404_),
    .ZN(_1405_));
 NOR2_X1 _2334_ (.A1(_1135_),
    .A2(_1314_),
    .ZN(_1406_));
 AOI21_X1 _2335_ (.A(_1406_),
    .B1(_1328_),
    .B2(_1135_),
    .ZN(_1407_));
 OAI21_X1 _2336_ (.A(_1405_),
    .B1(_1407_),
    .B2(_1384_),
    .ZN(_1408_));
 MUX2_X1 _2337_ (.A(_1389_),
    .B(_1401_),
    .S(_1408_),
    .Z(_1409_));
 NOR2_X1 _2338_ (.A1(_1400_),
    .A2(_1389_),
    .ZN(_1410_));
 AND2_X1 _2339_ (.A1(_1187_),
    .A2(_1219_),
    .ZN(_1411_));
 NAND3_X1 _2340_ (.A1(_1207_),
    .A2(_1379_),
    .A3(_1411_),
    .ZN(_1412_));
 OAI21_X1 _2341_ (.A(_1412_),
    .B1(_1411_),
    .B2(_1379_),
    .ZN(_1413_));
 AOI221_X2 _2342_ (.A(_1410_),
    .B1(_1202_),
    .B2(_1189_),
    .C1(_1947_),
    .C2(_1413_),
    .ZN(_1414_));
 NAND2_X1 _2343_ (.A1(_1409_),
    .A2(_1414_),
    .ZN(_1585_));
 NAND2_X1 _2344_ (.A1(net46),
    .A2(net91),
    .ZN(_1415_));
 XNOR2_X2 _2345_ (.A(_1222_),
    .B(_1415_),
    .ZN(_1896_));
 INV_X1 _2346_ (.A(_1896_),
    .ZN(_1586_));
 TAPCELL_X1 PHY_92 ();
 NAND3_X4 _2348_ (.A1(_1947_),
    .A2(_1187_),
    .A3(_1207_),
    .ZN(_1417_));
 NOR2_X1 _2349_ (.A1(_1355_),
    .A2(_1187_),
    .ZN(_1418_));
 AOI221_X1 _2350_ (.A(_1139_),
    .B1(_1187_),
    .B2(_1375_),
    .C1(_1418_),
    .C2(_1338_),
    .ZN(_1419_));
 TAPCELL_X1 PHY_91 ();
 TAPCELL_X1 PHY_90 ();
 MUX2_X1 _2353_ (.A(net45),
    .B(net44),
    .S(net94),
    .Z(_1422_));
 MUX2_X1 _2354_ (.A(_1396_),
    .B(_1422_),
    .S(_1135_),
    .Z(_1423_));
 NAND2_X1 _2355_ (.A1(_1365_),
    .A2(_1423_),
    .ZN(_1424_));
 OAI21_X1 _2356_ (.A(_1139_),
    .B1(_1205_),
    .B2(_1424_),
    .ZN(_1425_));
 AOI21_X1 _2357_ (.A(_1425_),
    .B1(_1418_),
    .B2(_1353_),
    .ZN(_1426_));
 OAI33_X1 _2358_ (.A1(_1185_),
    .A2(_1315_),
    .A3(_1417_),
    .B1(_1419_),
    .B2(_1426_),
    .B3(_1208_),
    .ZN(_1427_));
 XNOR2_X1 _2359_ (.A(_1379_),
    .B(_1427_),
    .ZN(_1591_));
 NAND2_X1 _2360_ (.A1(net44),
    .A2(net91),
    .ZN(_1428_));
 XNOR2_X1 _2361_ (.A(_1222_),
    .B(_1428_),
    .ZN(_1903_));
 INV_X1 _2362_ (.A(_1903_),
    .ZN(_1590_));
 NAND2_X1 _2363_ (.A1(_1134_),
    .A2(_1139_),
    .ZN(_1429_));
 NOR3_X1 _2364_ (.A1(_1355_),
    .A2(_1314_),
    .A3(_1429_),
    .ZN(_1430_));
 TAPCELL_X1 PHY_89 ();
 AOI21_X1 _2366_ (.A(_1139_),
    .B1(_1217_),
    .B2(_1842_),
    .ZN(_1432_));
 NOR3_X1 _2367_ (.A1(_1134_),
    .A2(_1355_),
    .A3(_1432_),
    .ZN(_1433_));
 OR2_X1 _2368_ (.A1(_1138_),
    .A2(_1328_),
    .ZN(_1434_));
 AOI21_X2 _2369_ (.A(_1430_),
    .B1(_1433_),
    .B2(_1434_),
    .ZN(_1435_));
 OAI21_X1 _2370_ (.A(_1403_),
    .B1(_1336_),
    .B2(_1135_),
    .ZN(_1436_));
 NOR3_X1 _2371_ (.A1(_1139_),
    .A2(_1355_),
    .A3(_1436_),
    .ZN(_1437_));
 TAPCELL_X1 PHY_88 ();
 NOR2_X1 _2373_ (.A1(_1138_),
    .A2(_1393_),
    .ZN(_1439_));
 NOR3_X1 _2374_ (.A1(_1187_),
    .A2(_1437_),
    .A3(_1439_),
    .ZN(_1440_));
 TAPCELL_X1 PHY_87 ();
 NAND2_X1 _2376_ (.A1(net94),
    .A2(net42),
    .ZN(_1442_));
 TAPCELL_X1 PHY_86 ();
 INV_X1 _2378_ (.A(net43),
    .ZN(_1444_));
 OAI21_X1 _2379_ (.A(_1442_),
    .B1(_1444_),
    .B2(net94),
    .ZN(_1445_));
 MUX2_X1 _2380_ (.A(_1422_),
    .B(_1445_),
    .S(_1135_),
    .Z(_1446_));
 NAND3_X1 _2381_ (.A1(_1139_),
    .A2(_1365_),
    .A3(_1446_),
    .ZN(_1447_));
 OAI21_X1 _2382_ (.A(_1447_),
    .B1(_1398_),
    .B2(_1139_),
    .ZN(_1448_));
 OAI21_X1 _2383_ (.A(_1190_),
    .B1(_1448_),
    .B2(_1205_),
    .ZN(_1449_));
 OAI22_X2 _2384_ (.A1(_1417_),
    .A2(_1435_),
    .B1(_1440_),
    .B2(_1449_),
    .ZN(_1450_));
 XNOR2_X1 _2385_ (.A(_1379_),
    .B(_1450_),
    .ZN(_1595_));
 NAND2_X1 _2386_ (.A1(net42),
    .A2(net91),
    .ZN(_1451_));
 XNOR2_X2 _2387_ (.A(_1222_),
    .B(_1451_),
    .ZN(_1911_));
 INV_X1 _2388_ (.A(_1911_),
    .ZN(_1594_));
 NOR2_X1 _2389_ (.A1(_1307_),
    .A2(_1376_),
    .ZN(_1452_));
 NOR3_X1 _2390_ (.A1(_1142_),
    .A2(_1205_),
    .A3(_1189_),
    .ZN(_1453_));
 NOR2_X1 _2391_ (.A1(_1444_),
    .A2(_1135_),
    .ZN(_1454_));
 TAPCELL_X1 PHY_85 ();
 AOI21_X1 _2393_ (.A(_1454_),
    .B1(_1135_),
    .B2(net39),
    .ZN(_1456_));
 NOR2_X1 _2394_ (.A1(net94),
    .A2(_1456_),
    .ZN(_1457_));
 TAPCELL_X1 PHY_84 ();
 MUX2_X1 _2396_ (.A(net42),
    .B(net28),
    .S(_1135_),
    .Z(_1459_));
 AOI21_X1 _2397_ (.A(_1457_),
    .B1(_1459_),
    .B2(net94),
    .ZN(_1460_));
 NAND2_X1 _2398_ (.A1(_1139_),
    .A2(_1365_),
    .ZN(_1461_));
 OAI22_X2 _2399_ (.A1(_1139_),
    .A2(_1424_),
    .B1(_1460_),
    .B2(_1461_),
    .ZN(_1462_));
 AOI221_X2 _2400_ (.A(_1452_),
    .B1(_1453_),
    .B2(_1385_),
    .C1(_1209_),
    .C2(_1462_),
    .ZN(_1463_));
 XNOR2_X1 _2401_ (.A(_1202_),
    .B(_1463_),
    .ZN(_1600_));
 NAND2_X1 _2402_ (.A1(net28),
    .A2(net91),
    .ZN(_1464_));
 XNOR2_X2 _2403_ (.A(_1222_),
    .B(_1464_),
    .ZN(_1919_));
 INV_X1 _2404_ (.A(_1919_),
    .ZN(_1599_));
 INV_X1 _2405_ (.A(_1935_),
    .ZN(_1943_));
 AOI21_X1 _2406_ (.A(_1187_),
    .B1(_1139_),
    .B2(_1943_),
    .ZN(_1946_));
 INV_X1 _2407_ (.A(_1925_),
    .ZN(_1465_));
 AOI21_X1 _2408_ (.A(_1927_),
    .B1(_1928_),
    .B2(_1604_),
    .ZN(_1466_));
 INV_X1 _2409_ (.A(_1926_),
    .ZN(_1467_));
 OAI21_X1 _2410_ (.A(_1465_),
    .B1(_1466_),
    .B2(_1467_),
    .ZN(_1468_));
 INV_X1 _2411_ (.A(_1468_),
    .ZN(_1601_));
 TAPCELL_X1 PHY_83 ();
 INV_X1 _2413_ (.A(_1910_),
    .ZN(_1470_));
 INV_X1 _2414_ (.A(_1917_),
    .ZN(_1471_));
 AOI21_X1 _2415_ (.A(_1921_),
    .B1(_1468_),
    .B2(_1922_),
    .ZN(_1472_));
 INV_X1 _2416_ (.A(_1918_),
    .ZN(_1473_));
 OAI21_X1 _2417_ (.A(_1471_),
    .B1(_1472_),
    .B2(_1473_),
    .ZN(_1474_));
 AOI21_X2 _2418_ (.A(_1913_),
    .B1(_1474_),
    .B2(_1914_),
    .ZN(_1475_));
 NOR2_X1 _2419_ (.A1(_1470_),
    .A2(_1475_),
    .ZN(_1476_));
 NOR2_X1 _2420_ (.A1(_1909_),
    .A2(_1476_),
    .ZN(_1589_));
 TAPCELL_X1 PHY_82 ();
 AND2_X1 _2422_ (.A1(_1906_),
    .A2(_1909_),
    .ZN(_1478_));
 OAI21_X1 _2423_ (.A(_1902_),
    .B1(_1905_),
    .B2(_1478_),
    .ZN(_1479_));
 NOR3_X1 _2424_ (.A1(_1893_),
    .A2(_1897_),
    .A3(_1901_),
    .ZN(_1480_));
 NAND3_X1 _2425_ (.A1(_1902_),
    .A2(_1906_),
    .A3(_1910_),
    .ZN(_1481_));
 OAI211_X2 _2426_ (.A(_1479_),
    .B(_1480_),
    .C1(_1475_),
    .C2(_1481_),
    .ZN(_1482_));
 NOR3_X1 _2427_ (.A1(_1898_),
    .A2(_1893_),
    .A3(_1897_),
    .ZN(_1483_));
 NOR2_X1 _2428_ (.A1(_1894_),
    .A2(_1893_),
    .ZN(_1484_));
 NOR2_X1 _2429_ (.A1(_1483_),
    .A2(_1484_),
    .ZN(_1485_));
 NAND2_X1 _2430_ (.A1(_1482_),
    .A2(_1485_),
    .ZN(_1579_));
 TAPCELL_X1 PHY_81 ();
 NAND3_X1 _2432_ (.A1(_1882_),
    .A2(_1886_),
    .A3(_1890_),
    .ZN(_1487_));
 AOI21_X1 _2433_ (.A(_1885_),
    .B1(_1889_),
    .B2(_1886_),
    .ZN(_1488_));
 INV_X1 _2434_ (.A(_1882_),
    .ZN(_1489_));
 OAI22_X2 _2435_ (.A1(_1579_),
    .A2(_1487_),
    .B1(_1488_),
    .B2(_1489_),
    .ZN(_1490_));
 OR2_X1 _2436_ (.A1(_1881_),
    .A2(_1490_),
    .ZN(_1491_));
 TAPCELL_X1 PHY_80 ();
 AOI21_X1 _2438_ (.A(_1879_),
    .B1(_1491_),
    .B2(_1880_),
    .ZN(_1569_));
 TAPCELL_X1 PHY_79 ();
 AOI21_X1 _2440_ (.A(_1853_),
    .B1(_1855_),
    .B2(_1854_),
    .ZN(_1494_));
 NAND2_X1 _2441_ (.A1(_1854_),
    .A2(_1856_),
    .ZN(_1495_));
 OR3_X1 _2442_ (.A1(_1862_),
    .A2(_1859_),
    .A3(_1861_),
    .ZN(_1496_));
 OR3_X1 _2443_ (.A1(_1859_),
    .A2(_1861_),
    .A3(_1865_),
    .ZN(_1497_));
 TAPCELL_X1 PHY_78 ();
 NAND2_X1 _2445_ (.A1(_1866_),
    .A2(_1867_),
    .ZN(_1499_));
 NAND3_X1 _2446_ (.A1(_1866_),
    .A2(_1868_),
    .A3(_1872_),
    .ZN(_1500_));
 OR3_X1 _2447_ (.A1(_1880_),
    .A2(_1875_),
    .A3(_1879_),
    .ZN(_1501_));
 OR3_X1 _2448_ (.A1(_1875_),
    .A2(_1879_),
    .A3(_1881_),
    .ZN(_1502_));
 OAI221_X2 _2449_ (.A(_1501_),
    .B1(_1502_),
    .B2(_1490_),
    .C1(_1876_),
    .C2(_1875_),
    .ZN(_1503_));
 INV_X1 _2450_ (.A(_1871_),
    .ZN(_1504_));
 NAND2_X1 _2451_ (.A1(_1866_),
    .A2(_1868_),
    .ZN(_1505_));
 OAI221_X2 _2452_ (.A(_1499_),
    .B1(_1500_),
    .B2(_1503_),
    .C1(_1504_),
    .C2(_1505_),
    .ZN(_1506_));
 OAI221_X2 _2453_ (.A(_1496_),
    .B1(_1497_),
    .B2(_1506_),
    .C1(_1860_),
    .C2(_1859_),
    .ZN(_1507_));
 OAI21_X1 _2454_ (.A(_1494_),
    .B1(_1495_),
    .B2(_1507_),
    .ZN(_1549_));
 AOI21_X1 _2455_ (.A(_1849_),
    .B1(_1549_),
    .B2(_1850_),
    .ZN(_1508_));
 INV_X1 _2456_ (.A(_1508_),
    .ZN(_1509_));
 AOI21_X1 _2457_ (.A(_1847_),
    .B1(_1509_),
    .B2(_1848_),
    .ZN(_1544_));
 OAI21_X1 _2458_ (.A(_1479_),
    .B1(_1481_),
    .B2(_1475_),
    .ZN(_0000_));
 NOR2_X1 _2459_ (.A1(_1901_),
    .A2(_0000_),
    .ZN(_1584_));
 INV_X1 _2460_ (.A(_1474_),
    .ZN(_1596_));
 NOR2_X2 _2461_ (.A1(_1547_),
    .A2(_1613_),
    .ZN(_0001_));
 TAPCELL_X1 PHY_77 ();
 TAPCELL_X1 PHY_76 ();
 AND2_X1 _2464_ (.A1(_1548_),
    .A2(_1553_),
    .ZN(_0004_));
 XNOR2_X2 _2465_ (.A(_1557_),
    .B(_1854_),
    .ZN(_0005_));
 XNOR2_X2 _2466_ (.A(_1562_),
    .B(_1860_),
    .ZN(_0006_));
 TAPCELL_X1 PHY_75 ();
 INV_X1 _2468_ (.A(_1558_),
    .ZN(_0008_));
 OAI21_X1 _2469_ (.A(_0005_),
    .B1(_0006_),
    .B2(_0008_),
    .ZN(_0009_));
 XOR2_X2 _2470_ (.A(_1552_),
    .B(_1848_),
    .Z(_0010_));
 AOI221_X1 _2471_ (.A(_0001_),
    .B1(_0004_),
    .B2(_0009_),
    .C1(_0010_),
    .C2(_1548_),
    .ZN(_0011_));
 TAPCELL_X1 PHY_74 ();
 NAND4_X4 _2473_ (.A1(_1558_),
    .A2(_1563_),
    .A3(_0005_),
    .A4(_0006_),
    .ZN(_0013_));
 XNOR2_X2 _2474_ (.A(_1552_),
    .B(_1848_),
    .ZN(_0014_));
 OAI211_X4 _2475_ (.A(_0014_),
    .B(_0004_),
    .C1(_1547_),
    .C2(_1613_),
    .ZN(_0015_));
 TAPCELL_X1 PHY_73 ();
 XOR2_X2 _2477_ (.A(_1567_),
    .B(_1866_),
    .Z(_0017_));
 NOR2_X1 _2478_ (.A1(_1568_),
    .A2(_0017_),
    .ZN(_0018_));
 OR3_X1 _2479_ (.A1(_0013_),
    .A2(_0015_),
    .A3(_0018_),
    .ZN(_0019_));
 XNOR2_X2 _2480_ (.A(_1567_),
    .B(_1866_),
    .ZN(_0020_));
 XOR2_X2 _2481_ (.A(_1572_),
    .B(_1872_),
    .Z(_0021_));
 NAND2_X1 _2482_ (.A1(_0020_),
    .A2(_0021_),
    .ZN(_0022_));
 TAPCELL_X1 PHY_72 ();
 INV_X1 _2484_ (.A(_1573_),
    .ZN(_0024_));
 TAPCELL_X1 PHY_71 ();
 INV_X1 _2486_ (.A(_1578_),
    .ZN(_0026_));
 XNOR2_X2 _2487_ (.A(_1577_),
    .B(_1880_),
    .ZN(_0027_));
 AOI21_X1 _2488_ (.A(_0024_),
    .B1(_0026_),
    .B2(_0027_),
    .ZN(_0028_));
 INV_X1 _2489_ (.A(_1583_),
    .ZN(_0029_));
 XOR2_X2 _2490_ (.A(_1582_),
    .B(_1886_),
    .Z(_0030_));
 NAND3_X1 _2491_ (.A1(_0029_),
    .A2(_0027_),
    .A3(_0030_),
    .ZN(_0031_));
 AOI21_X1 _2492_ (.A(_0022_),
    .B1(_0028_),
    .B2(_0031_),
    .ZN(_0032_));
 OAI21_X1 _2493_ (.A(_0011_),
    .B1(_0019_),
    .B2(_0032_),
    .ZN(_0033_));
 TAPCELL_X1 PHY_70 ();
 INV_X1 _2495_ (.A(_1608_),
    .ZN(_0035_));
 TAPCELL_X1 PHY_69 ();
 TAPCELL_X1 PHY_68 ();
 NOR2_X1 _2498_ (.A1(_1611_),
    .A2(_1614_),
    .ZN(_0038_));
 XNOR2_X2 _2499_ (.A(_1607_),
    .B(_1926_),
    .ZN(_0039_));
 AND3_X1 _2500_ (.A1(_0035_),
    .A2(_0038_),
    .A3(_0039_),
    .ZN(_0040_));
 TAPCELL_X1 PHY_67 ();
 NAND2_X1 _2502_ (.A1(_1598_),
    .A2(_1603_),
    .ZN(_0042_));
 XNOR2_X2 _2503_ (.A(_1602_),
    .B(_1918_),
    .ZN(_0043_));
 XNOR2_X2 _2504_ (.A(_1597_),
    .B(_1910_),
    .ZN(_0044_));
 NOR3_X2 _2505_ (.A1(_0042_),
    .A2(_0043_),
    .A3(_0044_),
    .ZN(_0045_));
 TAPCELL_X1 PHY_66 ();
 TAPCELL_X1 PHY_65 ();
 XOR2_X2 _2508_ (.A(_1587_),
    .B(_1894_),
    .Z(_0048_));
 XOR2_X2 _2509_ (.A(_1592_),
    .B(_1902_),
    .Z(_0049_));
 AND4_X1 _2510_ (.A1(_1588_),
    .A2(_1593_),
    .A3(_0048_),
    .A4(_0049_),
    .ZN(_0050_));
 NAND3_X1 _2511_ (.A1(_0040_),
    .A2(_0045_),
    .A3(_0050_),
    .ZN(_0051_));
 NAND4_X4 _2512_ (.A1(_1583_),
    .A2(_1578_),
    .A3(_0027_),
    .A4(_0030_),
    .ZN(_0052_));
 NAND4_X4 _2513_ (.A1(_1573_),
    .A2(_1568_),
    .A3(_0020_),
    .A4(_0021_),
    .ZN(_0053_));
 NOR4_X4 _2514_ (.A1(_0013_),
    .A2(_0015_),
    .A3(_0052_),
    .A4(_0053_),
    .ZN(_0054_));
 NAND2_X2 _2515_ (.A1(_0051_),
    .A2(_0054_),
    .ZN(_1637_));
 XOR2_X2 _2516_ (.A(_1597_),
    .B(_1910_),
    .Z(_0055_));
 NAND2_X1 _2517_ (.A1(_0055_),
    .A2(_0049_),
    .ZN(_0056_));
 INV_X1 _2518_ (.A(_1611_),
    .ZN(_0057_));
 OAI21_X1 _2519_ (.A(_0039_),
    .B1(_1608_),
    .B2(_0057_),
    .ZN(_0058_));
 INV_X1 _2520_ (.A(_0042_),
    .ZN(_0059_));
 AOI221_X2 _2521_ (.A(_0056_),
    .B1(_0058_),
    .B2(_0059_),
    .C1(_0043_),
    .C2(_1598_),
    .ZN(_0060_));
 XNOR2_X2 _2522_ (.A(_1592_),
    .B(_1902_),
    .ZN(_0061_));
 OAI21_X1 _2523_ (.A(_1588_),
    .B1(_1593_),
    .B2(_0061_),
    .ZN(_0062_));
 OAI21_X2 _2524_ (.A(_0048_),
    .B1(_0060_),
    .B2(_0062_),
    .ZN(_0063_));
 OAI21_X4 _2525_ (.A(_0033_),
    .B1(_1637_),
    .B2(_0063_),
    .ZN(_0064_));
 INV_X8 _2526_ (.A(_0064_),
    .ZN(_0065_));
 TAPCELL_X1 PHY_64 ();
 TAPCELL_X1 PHY_63 ();
 INV_X1 _2529_ (.A(net32),
    .ZN(_1840_));
 INV_X1 _2530_ (.A(net33),
    .ZN(_1514_));
 MUX2_X2 _2531_ (.A(_1514_),
    .B(_1511_),
    .S(_1131_),
    .Z(_1661_));
 INV_X1 _2532_ (.A(net34),
    .ZN(_1522_));
 NAND2_X1 _2533_ (.A1(net34),
    .A2(_1123_),
    .ZN(_0067_));
 OAI21_X2 _2534_ (.A(_0067_),
    .B1(_1123_),
    .B2(_1519_),
    .ZN(_1654_));
 INV_X1 _2535_ (.A(_1654_),
    .ZN(_1657_));
 INV_X1 _2536_ (.A(net35),
    .ZN(_1784_));
 MUX2_X2 _2537_ (.A(net35),
    .B(_1785_),
    .S(_1131_),
    .Z(_1646_));
 INV_X1 _2538_ (.A(_1646_),
    .ZN(_1650_));
 INV_X1 _2539_ (.A(net36),
    .ZN(_1526_));
 MUX2_X1 _2540_ (.A(_1526_),
    .B(_1531_),
    .S(_1131_),
    .Z(_1642_));
 INV_X1 _2541_ (.A(net37),
    .ZN(_1775_));
 MUX2_X2 _2542_ (.A(_1775_),
    .B(_1535_),
    .S(_1131_),
    .Z(_0068_));
 TAPCELL_X1 PHY_62 ();
 INV_X4 _2544_ (.A(_0068_),
    .ZN(_1633_));
 INV_X1 _2545_ (.A(net38),
    .ZN(_1539_));
 MUX2_X2 _2546_ (.A(net38),
    .B(_1540_),
    .S(_1131_),
    .Z(_1673_));
 INV_X1 _2547_ (.A(_1673_),
    .ZN(_1632_));
 MUX2_X2 _2548_ (.A(net6),
    .B(net40),
    .S(_1123_),
    .Z(_1718_));
 AND4_X1 _2549_ (.A1(_1558_),
    .A2(_1563_),
    .A3(_0005_),
    .A4(_0006_),
    .ZN(_0070_));
 XOR2_X2 _2550_ (.A(_1577_),
    .B(_1880_),
    .Z(_0071_));
 XNOR2_X1 _2551_ (.A(_1582_),
    .B(_1886_),
    .ZN(_0072_));
 NOR4_X1 _2552_ (.A1(_0029_),
    .A2(_0026_),
    .A3(_0071_),
    .A4(_0072_),
    .ZN(_0073_));
 NAND4_X1 _2553_ (.A1(_1588_),
    .A2(_1593_),
    .A3(_0048_),
    .A4(_0049_),
    .ZN(_0074_));
 OAI211_X2 _2554_ (.A(_0070_),
    .B(_0073_),
    .C1(_0074_),
    .C2(_0045_),
    .ZN(_0075_));
 AOI21_X2 _2555_ (.A(_0015_),
    .B1(_0053_),
    .B2(_0070_),
    .ZN(_0076_));
 NAND2_X4 _2556_ (.A1(_0075_),
    .A2(_0076_),
    .ZN(_1653_));
 INV_X1 _2557_ (.A(_1653_),
    .ZN(_1656_));
 INV_X1 _2558_ (.A(_1637_),
    .ZN(_1641_));
 INV_X1 _2559_ (.A(_1640_),
    .ZN(_1628_));
 TAPCELL_X1 PHY_61 ();
 TAPCELL_X1 PHY_60 ();
 NAND2_X1 _2562_ (.A1(_0045_),
    .A2(_0050_),
    .ZN(_0078_));
 NOR2_X1 _2563_ (.A1(_0040_),
    .A2(_0078_),
    .ZN(_0079_));
 NOR3_X1 _2564_ (.A1(_0052_),
    .A2(_0053_),
    .A3(_0079_),
    .ZN(_0080_));
 OR3_X2 _2565_ (.A1(_0013_),
    .A2(_0015_),
    .A3(_0080_),
    .ZN(_1645_));
 INV_X1 _2566_ (.A(_1645_),
    .ZN(_1649_));
 OAI21_X1 _2567_ (.A(_1548_),
    .B1(_1613_),
    .B2(_1547_),
    .ZN(_0081_));
 NAND2_X1 _2568_ (.A1(_1558_),
    .A2(_0005_),
    .ZN(_0082_));
 AND2_X1 _2569_ (.A1(_1553_),
    .A2(_0014_),
    .ZN(_0083_));
 AOI21_X1 _2570_ (.A(_0081_),
    .B1(_0082_),
    .B2(_0083_),
    .ZN(_0084_));
 NAND2_X1 _2571_ (.A1(_1588_),
    .A2(_0048_),
    .ZN(_0085_));
 XOR2_X1 _2572_ (.A(_1607_),
    .B(_1926_),
    .Z(_0086_));
 OR3_X1 _2573_ (.A1(_1608_),
    .A2(_0038_),
    .A3(_0086_),
    .ZN(_0087_));
 INV_X1 _2574_ (.A(_1593_),
    .ZN(_0088_));
 INV_X1 _2575_ (.A(_1603_),
    .ZN(_0089_));
 NOR4_X1 _2576_ (.A1(_0088_),
    .A2(_0089_),
    .A3(_0043_),
    .A4(_0061_),
    .ZN(_0090_));
 NAND2_X1 _2577_ (.A1(_1598_),
    .A2(_0055_),
    .ZN(_0091_));
 NOR2_X1 _2578_ (.A1(_0088_),
    .A2(_0061_),
    .ZN(_0092_));
 AOI221_X2 _2579_ (.A(_0085_),
    .B1(_0087_),
    .B2(_0090_),
    .C1(_0091_),
    .C2(_0092_),
    .ZN(_0093_));
 OR4_X1 _2580_ (.A1(_0013_),
    .A2(_0015_),
    .A3(_0052_),
    .A4(_0053_),
    .ZN(_0094_));
 NAND2_X1 _2581_ (.A1(_0070_),
    .A2(_0083_),
    .ZN(_0095_));
 AND2_X1 _2582_ (.A1(_1568_),
    .A2(_0020_),
    .ZN(_0096_));
 OAI211_X2 _2583_ (.A(_1573_),
    .B(_0021_),
    .C1(_0071_),
    .C2(_0026_),
    .ZN(_0097_));
 AND2_X1 _2584_ (.A1(_0096_),
    .A2(_0097_),
    .ZN(_0098_));
 OAI221_X2 _2585_ (.A(_0084_),
    .B1(_0093_),
    .B2(_0094_),
    .C1(_0095_),
    .C2(_0098_),
    .ZN(_0099_));
 INV_X2 _2586_ (.A(_0099_),
    .ZN(_1660_));
 AND2_X1 _2587_ (.A1(_1648_),
    .A2(_1640_),
    .ZN(_0100_));
 OAI21_X1 _2588_ (.A(_0100_),
    .B1(_1658_),
    .B2(_1624_),
    .ZN(_0101_));
 NOR2_X1 _2589_ (.A1(_1658_),
    .A2(_1662_),
    .ZN(_0102_));
 INV_X1 _2590_ (.A(_1667_),
    .ZN(_0103_));
 OAI21_X1 _2591_ (.A(_1663_),
    .B1(_0103_),
    .B2(_1668_),
    .ZN(_0104_));
 AOI21_X2 _2592_ (.A(_0101_),
    .B1(_0102_),
    .B2(_0104_),
    .ZN(_0105_));
 AOI21_X2 _2593_ (.A(_1643_),
    .B1(_1651_),
    .B2(_1640_),
    .ZN(_0106_));
 INV_X1 _2594_ (.A(_0106_),
    .ZN(_0107_));
 OAI21_X4 _2595_ (.A(_1716_),
    .B1(_0105_),
    .B2(_0107_),
    .ZN(_0108_));
 NOR2_X4 _2596_ (.A1(_1633_),
    .A2(_0108_),
    .ZN(_0109_));
 NOR2_X1 _2597_ (.A1(_0051_),
    .A2(_0094_),
    .ZN(_0110_));
 INV_X1 _2598_ (.A(_1716_),
    .ZN(_0111_));
 OR2_X1 _2599_ (.A1(_1658_),
    .A2(_1662_),
    .ZN(_0112_));
 INV_X1 _2600_ (.A(_1663_),
    .ZN(_1620_));
 INV_X1 _2601_ (.A(_1668_),
    .ZN(_0113_));
 AOI21_X1 _2602_ (.A(_1620_),
    .B1(_1667_),
    .B2(_0113_),
    .ZN(_0114_));
 OAI221_X2 _2603_ (.A(_0100_),
    .B1(_0112_),
    .B2(_0114_),
    .C1(_1624_),
    .C2(_1658_),
    .ZN(_0115_));
 AOI21_X4 _2604_ (.A(_0111_),
    .B1(_0115_),
    .B2(_0106_),
    .ZN(_0116_));
 AOI21_X4 _2605_ (.A(_0110_),
    .B1(_0116_),
    .B2(_0068_),
    .ZN(_0117_));
 TAPCELL_X1 PHY_59 ();
 INV_X2 _2607_ (.A(_1671_),
    .ZN(_0119_));
 OAI22_X4 _2608_ (.A1(_1653_),
    .A2(_0109_),
    .B1(_0117_),
    .B2(_0119_),
    .ZN(_0120_));
 INV_X8 _2609_ (.A(_0120_),
    .ZN(_0121_));
 TAPCELL_X1 PHY_58 ();
 TAPCELL_X1 PHY_57 ();
 TAPCELL_X1 PHY_56 ();
 AND3_X1 _2613_ (.A1(_0040_),
    .A2(_0045_),
    .A3(_0050_),
    .ZN(_0124_));
 NAND2_X2 _2614_ (.A1(_0124_),
    .A2(_0054_),
    .ZN(_0125_));
 OAI21_X4 _2615_ (.A(_0125_),
    .B1(_0108_),
    .B2(_1633_),
    .ZN(_0126_));
 TAPCELL_X1 PHY_55 ();
 INV_X1 _2617_ (.A(_1642_),
    .ZN(_1638_));
 AND3_X1 _2618_ (.A1(_1669_),
    .A2(_1654_),
    .A3(_1646_),
    .ZN(_1676_));
 AND3_X1 _2619_ (.A1(_1638_),
    .A2(_1633_),
    .A3(_1676_),
    .ZN(_1672_));
 NAND3_X1 _2620_ (.A1(_1719_),
    .A2(_0126_),
    .A3(_1672_),
    .ZN(_1699_));
 INV_X1 _2621_ (.A(_1699_),
    .ZN(_1703_));
 TAPCELL_X1 PHY_54 ();
 TAPCELL_X1 PHY_53 ();
 OAI22_X4 _2624_ (.A1(_0054_),
    .A2(_0109_),
    .B1(_0117_),
    .B2(_1678_),
    .ZN(_1691_));
 XNOR2_X2 _2625_ (.A(_1677_),
    .B(_1633_),
    .ZN(_0130_));
 TAPCELL_X1 PHY_52 ();
 TAPCELL_X1 PHY_51 ();
 NAND2_X2 _2628_ (.A1(_0068_),
    .A2(_0116_),
    .ZN(_0133_));
 AOI221_X2 _2629_ (.A(_0130_),
    .B1(_0125_),
    .B2(_0133_),
    .C1(_1689_),
    .C2(_1691_),
    .ZN(_1694_));
 XOR2_X1 _2630_ (.A(_1674_),
    .B(_1718_),
    .Z(_0134_));
 AND2_X1 _2631_ (.A1(_1675_),
    .A2(_0126_),
    .ZN(_1695_));
 NAND3_X1 _2632_ (.A1(_1694_),
    .A2(_0134_),
    .A3(_1695_),
    .ZN(_1698_));
 INV_X1 _2633_ (.A(_1698_),
    .ZN(_1702_));
 INV_X1 _2634_ (.A(_1697_),
    .ZN(_0135_));
 XNOR2_X1 _2635_ (.A(_1674_),
    .B(_1718_),
    .ZN(_0136_));
 OAI21_X2 _2636_ (.A(_1696_),
    .B1(_0117_),
    .B2(_0136_),
    .ZN(_0137_));
 TAPCELL_X1 PHY_50 ();
 OR3_X2 _2638_ (.A1(_1696_),
    .A2(_0117_),
    .A3(_0136_),
    .ZN(_0139_));
 AND3_X4 _2639_ (.A1(_0135_),
    .A2(_0137_),
    .A3(_0139_),
    .ZN(_0140_));
 TAPCELL_X1 PHY_49 ();
 TAPCELL_X1 PHY_48 ();
 TAPCELL_X1 PHY_47 ();
 INV_X2 _2643_ (.A(_1692_),
    .ZN(_0144_));
 XNOR2_X2 _2644_ (.A(_1677_),
    .B(_0068_),
    .ZN(_0145_));
 AOI21_X4 _2645_ (.A(_0144_),
    .B1(_0126_),
    .B2(_0145_),
    .ZN(_0146_));
 NOR3_X4 _2646_ (.A1(_1692_),
    .A2(_0117_),
    .A3(_0130_),
    .ZN(_0147_));
 NOR2_X4 _2647_ (.A1(_0146_),
    .A2(_0147_),
    .ZN(_0148_));
 TAPCELL_X1 PHY_46 ();
 TAPCELL_X1 PHY_45 ();
 INV_X4 _2650_ (.A(_1693_),
    .ZN(_0151_));
 TAPCELL_X1 PHY_44 ();
 INV_X4 _2652_ (.A(net85),
    .ZN(_0153_));
 NAND2_X2 _2653_ (.A1(_0151_),
    .A2(_0153_),
    .ZN(_0154_));
 TAPCELL_X1 PHY_43 ();
 TAPCELL_X1 PHY_42 ();
 TAPCELL_X1 PHY_41 ();
 NAND2_X1 _2657_ (.A1(_1614_),
    .A2(net82),
    .ZN(_0158_));
 TAPCELL_X1 PHY_40 ();
 TAPCELL_X1 PHY_39 ();
 MUX2_X2 _2660_ (.A(net87),
    .B(_0064_),
    .S(net86),
    .Z(_0161_));
 TAPCELL_X1 PHY_38 ();
 OAI21_X1 _2662_ (.A(_0121_),
    .B1(_0158_),
    .B2(_0161_),
    .ZN(_0163_));
 INV_X8 _2663_ (.A(net82),
    .ZN(_0164_));
 TAPCELL_X1 PHY_37 ();
 TAPCELL_X1 PHY_36 ();
 TAPCELL_X1 PHY_35 ();
 MUX2_X1 _2667_ (.A(_1603_),
    .B(_0039_),
    .S(net87),
    .Z(_0168_));
 NOR3_X2 _2668_ (.A1(_0164_),
    .A2(net86),
    .A3(_0168_),
    .ZN(_0169_));
 NAND2_X1 _2669_ (.A1(net82),
    .A2(_0086_),
    .ZN(_0170_));
 AOI21_X1 _2670_ (.A(_0170_),
    .B1(_0116_),
    .B2(_0068_),
    .ZN(_0171_));
 NAND2_X1 _2671_ (.A1(_0089_),
    .A2(net82),
    .ZN(_0172_));
 AOI21_X1 _2672_ (.A(_0172_),
    .B1(_0116_),
    .B2(_0068_),
    .ZN(_0173_));
 MUX2_X1 _2673_ (.A(_0171_),
    .B(_0173_),
    .S(_0065_),
    .Z(_0174_));
 OR2_X1 _2674_ (.A1(_0169_),
    .A2(_0174_),
    .ZN(_0175_));
 TAPCELL_X1 PHY_34 ();
 NOR2_X1 _2676_ (.A1(_1683_),
    .A2(_0119_),
    .ZN(_0177_));
 INV_X1 _2677_ (.A(_0177_),
    .ZN(_0178_));
 NAND2_X1 _2678_ (.A1(_1656_),
    .A2(_0099_),
    .ZN(_0179_));
 MUX2_X2 _2679_ (.A(_0178_),
    .B(_0179_),
    .S(_0117_),
    .Z(_0180_));
 TAPCELL_X1 PHY_33 ();
 TAPCELL_X1 PHY_32 ();
 TAPCELL_X1 PHY_31 ();
 MUX2_X1 _2683_ (.A(_1608_),
    .B(_1611_),
    .S(net87),
    .Z(_0184_));
 NAND3_X1 _2684_ (.A1(net82),
    .A2(_0126_),
    .A3(_0184_),
    .ZN(_0185_));
 NOR2_X1 _2685_ (.A1(_0057_),
    .A2(_0164_),
    .ZN(_0186_));
 OAI21_X1 _2686_ (.A(_0186_),
    .B1(_0108_),
    .B2(_1633_),
    .ZN(_0187_));
 NOR2_X1 _2687_ (.A1(_0035_),
    .A2(_0164_),
    .ZN(_0188_));
 OAI21_X1 _2688_ (.A(_0188_),
    .B1(_0108_),
    .B2(_1633_),
    .ZN(_0189_));
 MUX2_X1 _2689_ (.A(_0187_),
    .B(_0189_),
    .S(_0065_),
    .Z(_0190_));
 AOI21_X1 _2690_ (.A(_0121_),
    .B1(_0185_),
    .B2(_0190_),
    .ZN(_0191_));
 INV_X1 _2691_ (.A(_1683_),
    .ZN(_0192_));
 MUX2_X2 _2692_ (.A(_0192_),
    .B(_0099_),
    .S(_0117_),
    .Z(_0193_));
 TAPCELL_X1 PHY_30 ();
 TAPCELL_X1 PHY_29 ();
 OAI221_X2 _2695_ (.A(_0163_),
    .B1(_0175_),
    .B2(_0180_),
    .C1(_0191_),
    .C2(_0193_),
    .ZN(_0196_));
 NAND2_X1 _2696_ (.A1(_1653_),
    .A2(_0099_),
    .ZN(_0197_));
 NAND2_X1 _2697_ (.A1(_0192_),
    .A2(_0119_),
    .ZN(_0198_));
 MUX2_X2 _2698_ (.A(_0197_),
    .B(_0198_),
    .S(_0126_),
    .Z(_0199_));
 TAPCELL_X1 PHY_28 ();
 TAPCELL_X1 PHY_27 ();
 MUX2_X1 _2701_ (.A(_1573_),
    .B(_0027_),
    .S(_1681_),
    .Z(_0202_));
 NOR3_X2 _2702_ (.A1(_0164_),
    .A2(net86),
    .A3(_0202_),
    .ZN(_0203_));
 NAND2_X1 _2703_ (.A1(net82),
    .A2(_0071_),
    .ZN(_0204_));
 TAPCELL_X1 PHY_26 ();
 TAPCELL_X1 PHY_25 ();
 AOI21_X1 _2706_ (.A(_0204_),
    .B1(_0116_),
    .B2(_0068_),
    .ZN(_0207_));
 NAND2_X1 _2707_ (.A1(_0024_),
    .A2(net82),
    .ZN(_0208_));
 AOI21_X1 _2708_ (.A(_0208_),
    .B1(_0116_),
    .B2(_0068_),
    .ZN(_0209_));
 MUX2_X1 _2709_ (.A(_0207_),
    .B(_0209_),
    .S(_0065_),
    .Z(_0210_));
 NOR3_X1 _2710_ (.A1(_0199_),
    .A2(_0203_),
    .A3(_0210_),
    .ZN(_0211_));
 MUX2_X1 _2711_ (.A(_1568_),
    .B(_0021_),
    .S(_1681_),
    .Z(_0212_));
 NOR3_X2 _2712_ (.A1(_0164_),
    .A2(_0117_),
    .A3(_0212_),
    .ZN(_0213_));
 AOI211_X4 _2713_ (.A(_0164_),
    .B(_0021_),
    .C1(_0068_),
    .C2(_0116_),
    .ZN(_0214_));
 OR2_X1 _2714_ (.A1(_1568_),
    .A2(_0164_),
    .ZN(_0215_));
 AOI21_X1 _2715_ (.A(_0215_),
    .B1(_0116_),
    .B2(_0068_),
    .ZN(_0216_));
 MUX2_X1 _2716_ (.A(_0214_),
    .B(_0216_),
    .S(_0065_),
    .Z(_0217_));
 NOR4_X1 _2717_ (.A1(_0121_),
    .A2(_0193_),
    .A3(_0213_),
    .A4(_0217_),
    .ZN(_0218_));
 MUX2_X1 _2718_ (.A(_1563_),
    .B(_0020_),
    .S(_1681_),
    .Z(_0219_));
 NOR3_X2 _2719_ (.A1(_0164_),
    .A2(_0117_),
    .A3(_0219_),
    .ZN(_0220_));
 NAND2_X1 _2720_ (.A1(net82),
    .A2(_0017_),
    .ZN(_0221_));
 AOI21_X1 _2721_ (.A(_0221_),
    .B1(_0116_),
    .B2(_0068_),
    .ZN(_0222_));
 OR2_X1 _2722_ (.A1(_1563_),
    .A2(_0164_),
    .ZN(_0223_));
 AOI21_X1 _2723_ (.A(_0223_),
    .B1(_0116_),
    .B2(_0068_),
    .ZN(_0224_));
 MUX2_X1 _2724_ (.A(_0222_),
    .B(_0224_),
    .S(_0065_),
    .Z(_0225_));
 MUX2_X1 _2725_ (.A(_1578_),
    .B(_0030_),
    .S(_1681_),
    .Z(_0226_));
 NOR3_X2 _2726_ (.A1(_0164_),
    .A2(net86),
    .A3(_0226_),
    .ZN(_0227_));
 NAND2_X1 _2727_ (.A1(net82),
    .A2(_0072_),
    .ZN(_0228_));
 AOI21_X1 _2728_ (.A(_0228_),
    .B1(_0116_),
    .B2(_0068_),
    .ZN(_0229_));
 NAND2_X1 _2729_ (.A1(_0026_),
    .A2(net82),
    .ZN(_0230_));
 AOI21_X1 _2730_ (.A(_0230_),
    .B1(_0116_),
    .B2(_0068_),
    .ZN(_0231_));
 MUX2_X1 _2731_ (.A(_0229_),
    .B(_0231_),
    .S(_0065_),
    .Z(_0232_));
 NAND2_X1 _2732_ (.A1(_1683_),
    .A2(_0119_),
    .ZN(_0233_));
 NAND2_X1 _2733_ (.A1(_1653_),
    .A2(_1660_),
    .ZN(_0234_));
 MUX2_X2 _2734_ (.A(_0233_),
    .B(_0234_),
    .S(_0117_),
    .Z(_0235_));
 TAPCELL_X1 PHY_24 ();
 OAI33_X1 _2736_ (.A1(_0180_),
    .A2(_0220_),
    .A3(_0225_),
    .B1(_0227_),
    .B2(_0232_),
    .B3(_0235_),
    .ZN(_0237_));
 OR3_X2 _2737_ (.A1(_0211_),
    .A2(_0218_),
    .A3(_0237_),
    .ZN(_0238_));
 OR2_X1 _2738_ (.A1(_1588_),
    .A2(net87),
    .ZN(_0239_));
 OR2_X1 _2739_ (.A1(_1588_),
    .A2(_0164_),
    .ZN(_0240_));
 OAI33_X1 _2740_ (.A1(_0164_),
    .A2(net86),
    .A3(_0239_),
    .B1(_0240_),
    .B2(_0109_),
    .B3(_0064_),
    .ZN(_0241_));
 NAND2_X1 _2741_ (.A1(net87),
    .A2(net82),
    .ZN(_0242_));
 NAND2_X1 _2742_ (.A1(net82),
    .A2(_0061_),
    .ZN(_0243_));
 OAI33_X1 _2743_ (.A1(_0049_),
    .A2(net86),
    .A3(_0242_),
    .B1(_0243_),
    .B2(_0109_),
    .B3(_0065_),
    .ZN(_0244_));
 NOR4_X1 _2744_ (.A1(_0121_),
    .A2(_0193_),
    .A3(_0241_),
    .A4(_0244_),
    .ZN(_0245_));
 TAPCELL_X1 PHY_23 ();
 XOR2_X1 _2746_ (.A(_1602_),
    .B(_1918_),
    .Z(_0247_));
 MUX2_X1 _2747_ (.A(_1598_),
    .B(_0247_),
    .S(net87),
    .Z(_0248_));
 NOR3_X2 _2748_ (.A1(_0164_),
    .A2(net86),
    .A3(_0248_),
    .ZN(_0249_));
 NAND2_X1 _2749_ (.A1(net82),
    .A2(_0043_),
    .ZN(_0250_));
 AOI21_X1 _2750_ (.A(_0250_),
    .B1(_0116_),
    .B2(_0068_),
    .ZN(_0251_));
 INV_X1 _2751_ (.A(_1598_),
    .ZN(_0252_));
 NAND2_X1 _2752_ (.A1(_0252_),
    .A2(net82),
    .ZN(_0253_));
 AOI21_X1 _2753_ (.A(_0253_),
    .B1(_0116_),
    .B2(_0068_),
    .ZN(_0254_));
 MUX2_X1 _2754_ (.A(_0251_),
    .B(_0254_),
    .S(_0065_),
    .Z(_0255_));
 MUX2_X1 _2755_ (.A(_1593_),
    .B(_0055_),
    .S(net87),
    .Z(_0256_));
 NOR3_X2 _2756_ (.A1(_0164_),
    .A2(net86),
    .A3(_0256_),
    .ZN(_0257_));
 NAND2_X1 _2757_ (.A1(net82),
    .A2(_0044_),
    .ZN(_0258_));
 AOI21_X1 _2758_ (.A(_0258_),
    .B1(_0116_),
    .B2(_0068_),
    .ZN(_0259_));
 NAND2_X1 _2759_ (.A1(_0088_),
    .A2(net82),
    .ZN(_0260_));
 AOI21_X1 _2760_ (.A(_0260_),
    .B1(_0116_),
    .B2(_0068_),
    .ZN(_0261_));
 MUX2_X1 _2761_ (.A(_0259_),
    .B(_0261_),
    .S(_0065_),
    .Z(_0262_));
 OAI33_X1 _2762_ (.A1(_0235_),
    .A2(_0249_),
    .A3(_0255_),
    .B1(_0257_),
    .B2(_0262_),
    .B3(_0199_),
    .ZN(_0263_));
 MUX2_X1 _2763_ (.A(_1583_),
    .B(_0048_),
    .S(_1681_),
    .Z(_0264_));
 NOR3_X2 _2764_ (.A1(_0164_),
    .A2(net86),
    .A3(_0264_),
    .ZN(_0265_));
 XNOR2_X1 _2765_ (.A(_1587_),
    .B(_1894_),
    .ZN(_0266_));
 NAND2_X1 _2766_ (.A1(net82),
    .A2(_0266_),
    .ZN(_0267_));
 AOI21_X1 _2767_ (.A(_0267_),
    .B1(_0116_),
    .B2(_0068_),
    .ZN(_0268_));
 NAND2_X1 _2768_ (.A1(_0029_),
    .A2(net82),
    .ZN(_0269_));
 AOI21_X1 _2769_ (.A(_0269_),
    .B1(_0116_),
    .B2(_0068_),
    .ZN(_0270_));
 MUX2_X1 _2770_ (.A(_0268_),
    .B(_0270_),
    .S(_0065_),
    .Z(_0271_));
 NOR3_X1 _2771_ (.A1(_0180_),
    .A2(_0265_),
    .A3(_0271_),
    .ZN(_0272_));
 OR3_X2 _2772_ (.A1(_0245_),
    .A2(_0263_),
    .A3(_0272_),
    .ZN(_0273_));
 TAPCELL_X1 PHY_22 ();
 TAPCELL_X1 PHY_21 ();
 MUX2_X1 _2775_ (.A(_0238_),
    .B(_0273_),
    .S(net84),
    .Z(_0276_));
 TAPCELL_X1 PHY_20 ();
 OAI221_X1 _2777_ (.A(_0148_),
    .B1(_0154_),
    .B2(_0196_),
    .C1(_0276_),
    .C2(_0151_),
    .ZN(_0278_));
 OAI21_X2 _2778_ (.A(_1692_),
    .B1(_0117_),
    .B2(_0130_),
    .ZN(_0279_));
 NAND3_X2 _2779_ (.A1(_0144_),
    .A2(_0126_),
    .A3(_0145_),
    .ZN(_0280_));
 NAND2_X4 _2780_ (.A1(_0279_),
    .A2(_0280_),
    .ZN(_0281_));
 TAPCELL_X1 PHY_19 ();
 NAND2_X4 _2782_ (.A1(_0151_),
    .A2(net84),
    .ZN(_0283_));
 INV_X1 _2783_ (.A(_1548_),
    .ZN(_0284_));
 MUX2_X1 _2784_ (.A(_0284_),
    .B(_0010_),
    .S(_1681_),
    .Z(_0285_));
 NAND2_X1 _2785_ (.A1(_1683_),
    .A2(_0285_),
    .ZN(_0286_));
 NAND3_X1 _2786_ (.A1(_0192_),
    .A2(_1681_),
    .A3(_0001_),
    .ZN(_0287_));
 NAND2_X1 _2787_ (.A1(_0286_),
    .A2(_0287_),
    .ZN(_0288_));
 AND3_X1 _2788_ (.A1(_1700_),
    .A2(_0109_),
    .A3(_0288_),
    .ZN(_0289_));
 MUX2_X1 _2789_ (.A(_1553_),
    .B(_0005_),
    .S(_1681_),
    .Z(_0290_));
 NOR3_X1 _2790_ (.A1(_0164_),
    .A2(_0117_),
    .A3(_0290_),
    .ZN(_0291_));
 XOR2_X1 _2791_ (.A(_1557_),
    .B(_1854_),
    .Z(_0292_));
 NAND2_X1 _2792_ (.A1(net82),
    .A2(_0292_),
    .ZN(_0293_));
 AOI21_X1 _2793_ (.A(_0293_),
    .B1(_0116_),
    .B2(_0068_),
    .ZN(_0294_));
 OR2_X1 _2794_ (.A1(_1553_),
    .A2(_0164_),
    .ZN(_0295_));
 AOI21_X1 _2795_ (.A(_0295_),
    .B1(_0116_),
    .B2(_0068_),
    .ZN(_0296_));
 MUX2_X1 _2796_ (.A(_0294_),
    .B(_0296_),
    .S(_0065_),
    .Z(_0297_));
 OR2_X1 _2797_ (.A1(_0291_),
    .A2(_0297_),
    .ZN(_0298_));
 MUX2_X1 _2798_ (.A(_1558_),
    .B(_0006_),
    .S(_1681_),
    .Z(_0299_));
 NOR3_X2 _2799_ (.A1(_0164_),
    .A2(_0117_),
    .A3(_0299_),
    .ZN(_0300_));
 XOR2_X1 _2800_ (.A(_1562_),
    .B(_1860_),
    .Z(_0301_));
 NAND2_X1 _2801_ (.A1(net82),
    .A2(_0301_),
    .ZN(_0302_));
 AOI21_X1 _2802_ (.A(_0302_),
    .B1(_0116_),
    .B2(_0068_),
    .ZN(_0303_));
 NAND2_X1 _2803_ (.A1(_0008_),
    .A2(net82),
    .ZN(_0304_));
 AOI21_X1 _2804_ (.A(_0304_),
    .B1(_0116_),
    .B2(_0068_),
    .ZN(_0305_));
 MUX2_X1 _2805_ (.A(_0303_),
    .B(_0305_),
    .S(_0065_),
    .Z(_0306_));
 OR2_X1 _2806_ (.A1(_0300_),
    .A2(_0306_),
    .ZN(_0307_));
 OAI222_X2 _2807_ (.A1(_0121_),
    .A2(_0289_),
    .B1(_0199_),
    .B2(_0298_),
    .C1(_0235_),
    .C2(_0307_),
    .ZN(_0308_));
 OAI21_X1 _2808_ (.A(_0281_),
    .B1(_0283_),
    .B2(_0308_),
    .ZN(_0309_));
 AND3_X1 _2809_ (.A1(_0140_),
    .A2(_0278_),
    .A3(_0309_),
    .ZN(_1760_));
 NAND3_X4 _2810_ (.A1(_0135_),
    .A2(_0137_),
    .A3(_0139_),
    .ZN(_0310_));
 TAPCELL_X1 PHY_18 ();
 NOR4_X1 _2812_ (.A1(_0121_),
    .A2(_0193_),
    .A3(_0291_),
    .A4(_0297_),
    .ZN(_0312_));
 NOR3_X1 _2813_ (.A1(_0235_),
    .A2(_0220_),
    .A3(_0225_),
    .ZN(_0313_));
 AND3_X1 _2814_ (.A1(_1700_),
    .A2(_0126_),
    .A3(_0285_),
    .ZN(_0314_));
 NAND2_X1 _2815_ (.A1(_1700_),
    .A2(_0010_),
    .ZN(_0315_));
 AOI21_X1 _2816_ (.A(_0315_),
    .B1(_0116_),
    .B2(_0068_),
    .ZN(_0316_));
 NAND2_X1 _2817_ (.A1(_0284_),
    .A2(_1700_),
    .ZN(_0317_));
 AOI21_X1 _2818_ (.A(_0317_),
    .B1(_0116_),
    .B2(_0068_),
    .ZN(_0318_));
 MUX2_X1 _2819_ (.A(_0316_),
    .B(_0318_),
    .S(_0065_),
    .Z(_0319_));
 OAI33_X1 _2820_ (.A1(_0199_),
    .A2(_0300_),
    .A3(_0306_),
    .B1(_0180_),
    .B2(_0314_),
    .B3(_0319_),
    .ZN(_0320_));
 OR4_X1 _2821_ (.A1(_0153_),
    .A2(_0312_),
    .A3(_0313_),
    .A4(_0320_),
    .ZN(_0321_));
 NAND2_X1 _2822_ (.A1(_1700_),
    .A2(_0001_),
    .ZN(_0322_));
 NOR3_X1 _2823_ (.A1(_1687_),
    .A2(_0322_),
    .A3(_0235_),
    .ZN(_0323_));
 AOI21_X1 _2824_ (.A(_0148_),
    .B1(_0161_),
    .B2(_0323_),
    .ZN(_0324_));
 NAND2_X1 _2825_ (.A1(_0321_),
    .A2(_0324_),
    .ZN(_0325_));
 TAPCELL_X1 PHY_17 ();
 NOR2_X1 _2827_ (.A1(_1687_),
    .A2(_0121_),
    .ZN(_0327_));
 NOR3_X1 _2828_ (.A1(_0193_),
    .A2(_0158_),
    .A3(_0161_),
    .ZN(_0328_));
 MUX2_X2 _2829_ (.A(_1683_),
    .B(_1660_),
    .S(net86),
    .Z(_0329_));
 AOI21_X1 _2830_ (.A(_0329_),
    .B1(_0185_),
    .B2(_0190_),
    .ZN(_0330_));
 OAI21_X1 _2831_ (.A(_0327_),
    .B1(_0328_),
    .B2(_0330_),
    .ZN(_0331_));
 AOI21_X1 _2832_ (.A(_1693_),
    .B1(_0148_),
    .B2(_0331_),
    .ZN(_0332_));
 NOR4_X1 _2833_ (.A1(_0121_),
    .A2(_0193_),
    .A3(_0203_),
    .A4(_0210_),
    .ZN(_0333_));
 NOR3_X1 _2834_ (.A1(_0235_),
    .A2(_0265_),
    .A3(_0271_),
    .ZN(_0334_));
 OAI33_X1 _2835_ (.A1(_0213_),
    .A2(_0217_),
    .A3(_0180_),
    .B1(_0227_),
    .B2(_0232_),
    .B3(_0199_),
    .ZN(_0335_));
 OR3_X1 _2836_ (.A1(_0333_),
    .A2(_0334_),
    .A3(_0335_),
    .ZN(_0336_));
 OR2_X1 _2837_ (.A1(_1687_),
    .A2(_0336_),
    .ZN(_0337_));
 NOR3_X1 _2838_ (.A1(_0235_),
    .A2(_0169_),
    .A3(_0174_),
    .ZN(_0338_));
 NOR4_X1 _2839_ (.A1(_0121_),
    .A2(_0193_),
    .A3(_0257_),
    .A4(_0262_),
    .ZN(_0339_));
 OAI33_X1 _2840_ (.A1(_0180_),
    .A2(_0241_),
    .A3(_0244_),
    .B1(_0249_),
    .B2(_0255_),
    .B3(_0199_),
    .ZN(_0340_));
 OR3_X1 _2841_ (.A1(_0338_),
    .A2(_0339_),
    .A3(_0340_),
    .ZN(_0341_));
 TAPCELL_X1 PHY_16 ();
 OAI21_X1 _2843_ (.A(_0337_),
    .B1(_0341_),
    .B2(_0153_),
    .ZN(_0343_));
 NOR3_X2 _2844_ (.A1(_0151_),
    .A2(_0146_),
    .A3(_0147_),
    .ZN(_0344_));
 AOI22_X2 _2845_ (.A1(_0325_),
    .A2(_0332_),
    .B1(_0343_),
    .B2(_0344_),
    .ZN(_0345_));
 NOR2_X1 _2846_ (.A1(_0310_),
    .A2(_0345_),
    .ZN(_1756_));
 NOR2_X2 _2847_ (.A1(_1693_),
    .A2(net85),
    .ZN(_0346_));
 NOR4_X1 _2848_ (.A1(_1692_),
    .A2(_1671_),
    .A3(_0117_),
    .A4(_0130_),
    .ZN(_0347_));
 AOI21_X1 _2849_ (.A(_1653_),
    .B1(_0116_),
    .B2(_0068_),
    .ZN(_0348_));
 NAND2_X1 _2850_ (.A1(_1692_),
    .A2(_0119_),
    .ZN(_0349_));
 OAI33_X1 _2851_ (.A1(_0144_),
    .A2(_1656_),
    .A3(_0126_),
    .B1(_0348_),
    .B2(_0145_),
    .B3(_0349_),
    .ZN(_0350_));
 OAI21_X1 _2852_ (.A(_0289_),
    .B1(_0347_),
    .B2(_0350_),
    .ZN(_0351_));
 NOR2_X1 _2853_ (.A1(_1653_),
    .A2(_1660_),
    .ZN(_0352_));
 MUX2_X2 _2854_ (.A(_0177_),
    .B(_0352_),
    .S(_0117_),
    .Z(_0353_));
 AND2_X1 _2855_ (.A1(_1614_),
    .A2(net82),
    .ZN(_0354_));
 INV_X4 _2856_ (.A(net87),
    .ZN(_0355_));
 TAPCELL_X1 PHY_15 ();
 MUX2_X2 _2858_ (.A(_0355_),
    .B(_0065_),
    .S(net86),
    .Z(_0357_));
 TAPCELL_X1 PHY_14 ();
 NAND3_X2 _2860_ (.A1(_0353_),
    .A2(_0354_),
    .A3(_0357_),
    .ZN(_0359_));
 OAI21_X1 _2861_ (.A(_0351_),
    .B1(_0359_),
    .B2(_0281_),
    .ZN(_0360_));
 NOR2_X1 _2862_ (.A1(_0148_),
    .A2(_0283_),
    .ZN(_0361_));
 OAI33_X1 _2863_ (.A1(_0235_),
    .A2(_0213_),
    .A3(_0217_),
    .B1(_0220_),
    .B2(_0225_),
    .B3(_0199_),
    .ZN(_0362_));
 NOR2_X4 _2864_ (.A1(_0121_),
    .A2(_0193_),
    .ZN(_0363_));
 NOR2_X1 _2865_ (.A1(_0300_),
    .A2(_0306_),
    .ZN(_0364_));
 NOR2_X1 _2866_ (.A1(_0291_),
    .A2(_0297_),
    .ZN(_0365_));
 AOI221_X2 _2867_ (.A(_0362_),
    .B1(_0363_),
    .B2(_0364_),
    .C1(_0365_),
    .C2(_0353_),
    .ZN(_0366_));
 AOI22_X1 _2868_ (.A1(_0346_),
    .A2(_0360_),
    .B1(_0361_),
    .B2(_0366_),
    .ZN(_0367_));
 NOR3_X1 _2869_ (.A1(_0203_),
    .A2(_0210_),
    .A3(_0180_),
    .ZN(_0368_));
 NOR4_X1 _2870_ (.A1(_0121_),
    .A2(_0193_),
    .A3(_0227_),
    .A4(_0232_),
    .ZN(_0369_));
 OAI33_X1 _2871_ (.A1(_0235_),
    .A2(_0241_),
    .A3(_0244_),
    .B1(_0265_),
    .B2(_0271_),
    .B3(_0199_),
    .ZN(_0370_));
 NOR2_X1 _2872_ (.A1(_0151_),
    .A2(net84),
    .ZN(_0371_));
 NAND3_X2 _2873_ (.A1(_0279_),
    .A2(_0280_),
    .A3(_0371_),
    .ZN(_0372_));
 NOR4_X1 _2874_ (.A1(_0368_),
    .A2(_0369_),
    .A3(_0370_),
    .A4(_0372_),
    .ZN(_0373_));
 NOR4_X1 _2875_ (.A1(_0121_),
    .A2(_0193_),
    .A3(_0249_),
    .A4(_0255_),
    .ZN(_0374_));
 NOR3_X1 _2876_ (.A1(_0180_),
    .A2(_0257_),
    .A3(_0262_),
    .ZN(_0375_));
 AND3_X1 _2877_ (.A1(net82),
    .A2(_0126_),
    .A3(_0184_),
    .ZN(_0376_));
 NAND2_X1 _2878_ (.A1(_1611_),
    .A2(net82),
    .ZN(_0377_));
 AOI21_X1 _2879_ (.A(_0377_),
    .B1(_0116_),
    .B2(_0068_),
    .ZN(_0378_));
 NAND2_X1 _2880_ (.A1(_1608_),
    .A2(net82),
    .ZN(_0379_));
 AOI21_X1 _2881_ (.A(_0379_),
    .B1(_0116_),
    .B2(_0068_),
    .ZN(_0380_));
 MUX2_X1 _2882_ (.A(_0378_),
    .B(_0380_),
    .S(_0065_),
    .Z(_0381_));
 OAI33_X1 _2883_ (.A1(_0199_),
    .A2(_0169_),
    .A3(_0174_),
    .B1(_0376_),
    .B2(_0381_),
    .B3(_0235_),
    .ZN(_0382_));
 NOR3_X1 _2884_ (.A1(_0374_),
    .A2(_0375_),
    .A3(_0382_),
    .ZN(_0383_));
 NAND2_X2 _2885_ (.A1(_1693_),
    .A2(net85),
    .ZN(_0384_));
 NOR2_X1 _2886_ (.A1(_0281_),
    .A2(_0384_),
    .ZN(_0385_));
 AOI21_X1 _2887_ (.A(_0373_),
    .B1(_0383_),
    .B2(_0385_),
    .ZN(_0386_));
 AOI21_X1 _2888_ (.A(_0310_),
    .B1(_0367_),
    .B2(_0386_),
    .ZN(_1752_));
 OAI33_X1 _2889_ (.A1(_0180_),
    .A2(_0227_),
    .A3(_0232_),
    .B1(_0241_),
    .B2(_0244_),
    .B3(_0199_),
    .ZN(_0387_));
 NOR2_X1 _2890_ (.A1(_0265_),
    .A2(_0271_),
    .ZN(_0388_));
 NOR2_X1 _2891_ (.A1(_0192_),
    .A2(_1671_),
    .ZN(_0389_));
 NOR2_X1 _2892_ (.A1(_1656_),
    .A2(_0099_),
    .ZN(_0390_));
 MUX2_X2 _2893_ (.A(_0389_),
    .B(_0390_),
    .S(_0117_),
    .Z(_0391_));
 NOR2_X1 _2894_ (.A1(_0257_),
    .A2(_0262_),
    .ZN(_0392_));
 AOI221_X2 _2895_ (.A(_0387_),
    .B1(_0388_),
    .B2(_0363_),
    .C1(_0391_),
    .C2(_0392_),
    .ZN(_0393_));
 NOR2_X1 _2896_ (.A1(_0310_),
    .A2(_0372_),
    .ZN(_0394_));
 AND3_X1 _2897_ (.A1(net85),
    .A2(_0140_),
    .A3(_0344_),
    .ZN(_0395_));
 OAI33_X1 _2898_ (.A1(_0180_),
    .A2(_0249_),
    .A3(_0255_),
    .B1(_0376_),
    .B2(_0381_),
    .B3(_0199_),
    .ZN(_0396_));
 NOR2_X1 _2899_ (.A1(_0169_),
    .A2(_0174_),
    .ZN(_0397_));
 TAPCELL_X1 PHY_13 ();
 AOI21_X1 _2901_ (.A(_0120_),
    .B1(_0354_),
    .B2(_0357_),
    .ZN(_0398_));
 AOI221_X2 _2902_ (.A(_0396_),
    .B1(_0397_),
    .B2(_0363_),
    .C1(_0329_),
    .C2(_0398_),
    .ZN(_0399_));
 AOI22_X1 _2903_ (.A1(_0393_),
    .A2(_0394_),
    .B1(_0395_),
    .B2(_0399_),
    .ZN(_0400_));
 OAI33_X1 _2904_ (.A1(_0235_),
    .A2(_0203_),
    .A3(_0210_),
    .B1(_0180_),
    .B2(_0306_),
    .B3(_0300_),
    .ZN(_0401_));
 NOR3_X1 _2905_ (.A1(_0199_),
    .A2(_0213_),
    .A3(_0217_),
    .ZN(_0402_));
 NOR4_X1 _2906_ (.A1(_0121_),
    .A2(_0193_),
    .A3(_0220_),
    .A4(_0225_),
    .ZN(_0403_));
 OR3_X1 _2907_ (.A1(_0401_),
    .A2(_0402_),
    .A3(_0403_),
    .ZN(_0404_));
 NOR2_X2 _2908_ (.A1(net83),
    .A2(_0153_),
    .ZN(_0405_));
 NAND3_X2 _2909_ (.A1(_0140_),
    .A2(_0281_),
    .A3(_0405_),
    .ZN(_0406_));
 OAI21_X1 _2910_ (.A(_0346_),
    .B1(_0147_),
    .B2(_0146_),
    .ZN(_0407_));
 OR2_X2 _2911_ (.A1(_0310_),
    .A2(_0407_),
    .ZN(_0408_));
 OR4_X1 _2912_ (.A1(_0192_),
    .A2(_0355_),
    .A3(_0133_),
    .A4(_0322_),
    .ZN(_0409_));
 NAND2_X1 _2913_ (.A1(_0120_),
    .A2(_0409_),
    .ZN(_0410_));
 OR2_X1 _2914_ (.A1(_0314_),
    .A2(_0319_),
    .ZN(_0411_));
 OAI221_X2 _2915_ (.A(_0410_),
    .B1(_0235_),
    .B2(_0298_),
    .C1(_0199_),
    .C2(_0411_),
    .ZN(_0412_));
 OAI221_X2 _2916_ (.A(_0400_),
    .B1(_0404_),
    .B2(_0406_),
    .C1(_0408_),
    .C2(_0412_),
    .ZN(_1749_));
 OR2_X1 _2917_ (.A1(_0310_),
    .A2(_0372_),
    .ZN(_0413_));
 NOR2_X1 _2918_ (.A1(_0273_),
    .A2(_0413_),
    .ZN(_0414_));
 NAND3_X1 _2919_ (.A1(net84),
    .A2(_0140_),
    .A3(_0344_),
    .ZN(_0415_));
 NOR2_X1 _2920_ (.A1(_0196_),
    .A2(_0415_),
    .ZN(_0416_));
 OAI22_X1 _2921_ (.A1(_0308_),
    .A2(_0408_),
    .B1(_0406_),
    .B2(_0238_),
    .ZN(_0417_));
 OR3_X1 _2922_ (.A1(_0414_),
    .A2(_0416_),
    .A3(_0417_),
    .ZN(_1745_));
 OR4_X1 _2923_ (.A1(_0312_),
    .A2(_0313_),
    .A3(_0320_),
    .A4(_0407_),
    .ZN(_0418_));
 NOR2_X1 _2924_ (.A1(_0330_),
    .A2(_0328_),
    .ZN(_0419_));
 NOR2_X1 _2925_ (.A1(_0151_),
    .A2(_0153_),
    .ZN(_0420_));
 NAND3_X1 _2926_ (.A1(_0120_),
    .A2(_0148_),
    .A3(_0420_),
    .ZN(_0421_));
 OAI221_X1 _2927_ (.A(_0418_),
    .B1(_0372_),
    .B2(_0341_),
    .C1(_0419_),
    .C2(_0421_),
    .ZN(_0422_));
 NAND2_X1 _2928_ (.A1(_0121_),
    .A2(_0420_),
    .ZN(_0423_));
 OAI22_X1 _2929_ (.A1(_0283_),
    .A2(_0336_),
    .B1(_0409_),
    .B2(_0423_),
    .ZN(_0424_));
 AOI21_X1 _2930_ (.A(_0422_),
    .B1(_0424_),
    .B2(_0281_),
    .ZN(_0425_));
 NOR2_X1 _2931_ (.A1(_0310_),
    .A2(_0425_),
    .ZN(_1740_));
 OR3_X1 _2932_ (.A1(_0374_),
    .A2(_0375_),
    .A3(_0382_),
    .ZN(_0426_));
 NAND2_X2 _2933_ (.A1(net83),
    .A2(_0153_),
    .ZN(_0427_));
 NOR2_X1 _2934_ (.A1(_0426_),
    .A2(_0427_),
    .ZN(_0428_));
 OAI21_X1 _2935_ (.A(_0148_),
    .B1(_0359_),
    .B2(_0384_),
    .ZN(_0429_));
 OAI21_X1 _2936_ (.A(_0140_),
    .B1(_0428_),
    .B2(_0429_),
    .ZN(_0430_));
 OR3_X1 _2937_ (.A1(_0368_),
    .A2(_0369_),
    .A3(_0370_),
    .ZN(_0431_));
 NAND3_X1 _2938_ (.A1(_1700_),
    .A2(_0109_),
    .A3(_0288_),
    .ZN(_0432_));
 OAI221_X2 _2939_ (.A(_0281_),
    .B1(_0283_),
    .B2(_0431_),
    .C1(_0423_),
    .C2(_0432_),
    .ZN(_0433_));
 AOI21_X2 _2940_ (.A(_0433_),
    .B1(_0366_),
    .B2(_0346_),
    .ZN(_0434_));
 NOR2_X1 _2941_ (.A1(_0430_),
    .A2(_0434_),
    .ZN(_1737_));
 AOI21_X1 _2942_ (.A(_0281_),
    .B1(_0371_),
    .B2(_0399_),
    .ZN(_0435_));
 OR2_X1 _2943_ (.A1(_0310_),
    .A2(_0435_),
    .ZN(_0436_));
 OR2_X1 _2944_ (.A1(_0153_),
    .A2(_0412_),
    .ZN(_0437_));
 NOR4_X1 _2945_ (.A1(_1687_),
    .A2(_0401_),
    .A3(_0402_),
    .A4(_0403_),
    .ZN(_0438_));
 AOI21_X1 _2946_ (.A(_0438_),
    .B1(_0393_),
    .B2(_1687_),
    .ZN(_0439_));
 MUX2_X1 _2947_ (.A(_0437_),
    .B(_0439_),
    .S(_0151_),
    .Z(_0440_));
 AOI21_X1 _2948_ (.A(_0436_),
    .B1(_0440_),
    .B2(_0281_),
    .ZN(_1732_));
 OAI21_X2 _2949_ (.A(_0148_),
    .B1(_0196_),
    .B2(_0427_),
    .ZN(_0441_));
 OAI21_X1 _2950_ (.A(_0281_),
    .B1(_0283_),
    .B2(_0273_),
    .ZN(_0442_));
 OAI22_X2 _2951_ (.A1(_0238_),
    .A2(_0154_),
    .B1(_0384_),
    .B2(_0308_),
    .ZN(_0443_));
 OAI211_X4 _2952_ (.A(_0140_),
    .B(_0441_),
    .C1(_0442_),
    .C2(_0443_),
    .ZN(_0444_));
 INV_X1 _2953_ (.A(_0444_),
    .ZN(_1729_));
 NAND3_X1 _2954_ (.A1(_1693_),
    .A2(_0321_),
    .A3(_0324_),
    .ZN(_0445_));
 NOR4_X1 _2955_ (.A1(_0121_),
    .A2(_0310_),
    .A3(_0419_),
    .A4(_0427_),
    .ZN(_0446_));
 NOR2_X1 _2956_ (.A1(_0310_),
    .A2(_0148_),
    .ZN(_0447_));
 AOI22_X1 _2957_ (.A1(_0405_),
    .A2(_0341_),
    .B1(_0336_),
    .B2(_0346_),
    .ZN(_0448_));
 OAI221_X2 _2958_ (.A(_0445_),
    .B1(_0446_),
    .B2(_0447_),
    .C1(_0448_),
    .C2(_0148_),
    .ZN(_0449_));
 INV_X1 _2959_ (.A(_0449_),
    .ZN(_1725_));
 MUX2_X1 _2960_ (.A(_0035_),
    .B(_0039_),
    .S(_0355_),
    .Z(_0450_));
 NOR3_X2 _2961_ (.A1(_0164_),
    .A2(net86),
    .A3(_0450_),
    .ZN(_0451_));
 MUX2_X1 _2962_ (.A(_0171_),
    .B(_0380_),
    .S(_0064_),
    .Z(_0452_));
 MUX2_X1 _2963_ (.A(_1593_),
    .B(_0049_),
    .S(_0355_),
    .Z(_0453_));
 NOR3_X2 _2964_ (.A1(_0164_),
    .A2(net86),
    .A3(_0453_),
    .ZN(_0454_));
 AOI21_X1 _2965_ (.A(_0243_),
    .B1(_0116_),
    .B2(_0068_),
    .ZN(_0455_));
 MUX2_X1 _2966_ (.A(_0455_),
    .B(_0261_),
    .S(_0064_),
    .Z(_0456_));
 OAI33_X1 _2967_ (.A1(_0235_),
    .A2(_0451_),
    .A3(_0452_),
    .B1(_0454_),
    .B2(_0456_),
    .B3(_0180_),
    .ZN(_0457_));
 MUX2_X1 _2968_ (.A(_0251_),
    .B(_0173_),
    .S(_0064_),
    .Z(_0458_));
 NAND3_X1 _2969_ (.A1(_0355_),
    .A2(net82),
    .A3(_0043_),
    .ZN(_0459_));
 NAND3_X1 _2970_ (.A1(_0089_),
    .A2(net87),
    .A3(net82),
    .ZN(_0460_));
 AOI21_X2 _2971_ (.A(_0133_),
    .B1(_0459_),
    .B2(_0460_),
    .ZN(_0461_));
 NOR3_X1 _2972_ (.A1(_0199_),
    .A2(_0458_),
    .A3(_0461_),
    .ZN(_0462_));
 MUX2_X1 _2973_ (.A(_1598_),
    .B(_0055_),
    .S(_0355_),
    .Z(_0463_));
 NOR3_X2 _2974_ (.A1(_0164_),
    .A2(net86),
    .A3(_0463_),
    .ZN(_0464_));
 MUX2_X1 _2975_ (.A(_0254_),
    .B(_0259_),
    .S(_0065_),
    .Z(_0465_));
 NOR4_X1 _2976_ (.A1(_0121_),
    .A2(_0193_),
    .A3(_0464_),
    .A4(_0465_),
    .ZN(_0466_));
 OR3_X1 _2977_ (.A1(_0457_),
    .A2(_0462_),
    .A3(_0466_),
    .ZN(_0467_));
 MUX2_X1 _2978_ (.A(_1573_),
    .B(_0021_),
    .S(_0355_),
    .Z(_0468_));
 NOR3_X2 _2979_ (.A1(_0164_),
    .A2(net86),
    .A3(_0468_),
    .ZN(_0469_));
 MUX2_X1 _2980_ (.A(_0209_),
    .B(_0214_),
    .S(_0065_),
    .Z(_0470_));
 NOR3_X1 _2981_ (.A1(_0180_),
    .A2(_0469_),
    .A3(_0470_),
    .ZN(_0471_));
 MUX2_X1 _2982_ (.A(_1583_),
    .B(_0030_),
    .S(_0355_),
    .Z(_0472_));
 NOR3_X2 _2983_ (.A1(_0164_),
    .A2(net86),
    .A3(_0472_),
    .ZN(_0473_));
 MUX2_X1 _2984_ (.A(_0229_),
    .B(_0270_),
    .S(_0064_),
    .Z(_0474_));
 MUX2_X1 _2985_ (.A(_1588_),
    .B(_0048_),
    .S(_0355_),
    .Z(_0475_));
 NOR3_X2 _2986_ (.A1(_0164_),
    .A2(net86),
    .A3(_0475_),
    .ZN(_0476_));
 AOI21_X1 _2987_ (.A(_0240_),
    .B1(_0116_),
    .B2(_0068_),
    .ZN(_0477_));
 MUX2_X1 _2988_ (.A(_0477_),
    .B(_0268_),
    .S(_0065_),
    .Z(_0478_));
 OAI33_X1 _2989_ (.A1(_0199_),
    .A2(_0473_),
    .A3(_0474_),
    .B1(_0476_),
    .B2(_0478_),
    .B3(_0235_),
    .ZN(_0479_));
 MUX2_X1 _2990_ (.A(_1578_),
    .B(_0027_),
    .S(_0355_),
    .Z(_0480_));
 NOR3_X2 _2991_ (.A1(_0164_),
    .A2(net86),
    .A3(_0480_),
    .ZN(_0481_));
 MUX2_X1 _2992_ (.A(_0207_),
    .B(_0231_),
    .S(_0064_),
    .Z(_0482_));
 NOR4_X1 _2993_ (.A1(_0121_),
    .A2(_0193_),
    .A3(_0481_),
    .A4(_0482_),
    .ZN(_0483_));
 OR3_X1 _2994_ (.A1(_0471_),
    .A2(_0479_),
    .A3(_0483_),
    .ZN(_0484_));
 MUX2_X1 _2995_ (.A(_0467_),
    .B(_0484_),
    .S(_0153_),
    .Z(_0485_));
 MUX2_X1 _2996_ (.A(_1553_),
    .B(_0014_),
    .S(_0355_),
    .Z(_0486_));
 NOR3_X2 _2997_ (.A1(_0164_),
    .A2(net86),
    .A3(_0486_),
    .ZN(_0487_));
 MUX2_X1 _2998_ (.A(_0296_),
    .B(_0316_),
    .S(_0065_),
    .Z(_0488_));
 NOR3_X1 _2999_ (.A1(_0180_),
    .A2(_0487_),
    .A3(_0488_),
    .ZN(_0489_));
 MUX2_X1 _3000_ (.A(_1568_),
    .B(_0020_),
    .S(_0355_),
    .Z(_0490_));
 NOR3_X1 _3001_ (.A1(_0164_),
    .A2(net86),
    .A3(_0490_),
    .ZN(_0491_));
 MUX2_X1 _3002_ (.A(_0216_),
    .B(_0222_),
    .S(_0065_),
    .Z(_0492_));
 MUX2_X1 _3003_ (.A(_1563_),
    .B(_0006_),
    .S(_0355_),
    .Z(_0493_));
 NOR3_X1 _3004_ (.A1(_0164_),
    .A2(net86),
    .A3(_0493_),
    .ZN(_0494_));
 MUX2_X1 _3005_ (.A(_0303_),
    .B(_0224_),
    .S(_0064_),
    .Z(_0495_));
 OAI33_X1 _3006_ (.A1(_0235_),
    .A2(_0491_),
    .A3(_0492_),
    .B1(_0494_),
    .B2(_0495_),
    .B3(_0199_),
    .ZN(_0496_));
 MUX2_X1 _3007_ (.A(_1558_),
    .B(_0005_),
    .S(_0355_),
    .Z(_0497_));
 NOR3_X2 _3008_ (.A1(_0164_),
    .A2(_0117_),
    .A3(_0497_),
    .ZN(_0498_));
 MUX2_X1 _3009_ (.A(_0294_),
    .B(_0305_),
    .S(_0064_),
    .Z(_0499_));
 NOR4_X1 _3010_ (.A1(_0121_),
    .A2(_0193_),
    .A3(_0498_),
    .A4(_0499_),
    .ZN(_0500_));
 OR3_X2 _3011_ (.A1(_0489_),
    .A2(_0496_),
    .A3(_0500_),
    .ZN(_0501_));
 MUX2_X1 _3012_ (.A(_0284_),
    .B(_0001_),
    .S(_0355_),
    .Z(_0502_));
 NAND4_X1 _3013_ (.A1(_1683_),
    .A2(_1700_),
    .A3(_0126_),
    .A4(_0502_),
    .ZN(_0503_));
 NOR2_X1 _3014_ (.A1(_0120_),
    .A2(_0503_),
    .ZN(_0504_));
 INV_X1 _3015_ (.A(_0504_),
    .ZN(_0505_));
 MUX2_X1 _3016_ (.A(_0501_),
    .B(_0505_),
    .S(_0153_),
    .Z(_0506_));
 MUX2_X1 _3017_ (.A(_0485_),
    .B(_0506_),
    .S(net83),
    .Z(_0507_));
 MUX2_X1 _3018_ (.A(_1611_),
    .B(_1614_),
    .S(net87),
    .Z(_0508_));
 NAND3_X1 _3019_ (.A1(net82),
    .A2(_0126_),
    .A3(_0508_),
    .ZN(_0509_));
 OAI21_X1 _3020_ (.A(_0354_),
    .B1(_0108_),
    .B2(_1633_),
    .ZN(_0510_));
 MUX2_X1 _3021_ (.A(_0510_),
    .B(_0187_),
    .S(_0065_),
    .Z(_0511_));
 NAND2_X1 _3022_ (.A1(_0509_),
    .A2(_0511_),
    .ZN(_0512_));
 NAND2_X1 _3023_ (.A1(_0353_),
    .A2(_0512_),
    .ZN(_0513_));
 OAI22_X1 _3024_ (.A1(_0148_),
    .A2(_0507_),
    .B1(_0513_),
    .B2(_0372_),
    .ZN(_0514_));
 AND2_X1 _3025_ (.A1(_0140_),
    .A2(_0514_),
    .ZN(_1722_));
 XOR2_X1 _3026_ (.A(_1626_),
    .B(_1709_),
    .Z(net67));
 AOI21_X1 _3027_ (.A(_1706_),
    .B1(_1707_),
    .B2(_1622_),
    .ZN(_0515_));
 INV_X1 _3028_ (.A(_0515_),
    .ZN(_0516_));
 AOI21_X1 _3029_ (.A(_1708_),
    .B1(_0516_),
    .B2(_1709_),
    .ZN(_1629_));
 XNOR2_X1 _3030_ (.A(_1631_),
    .B(_1714_),
    .ZN(net69));
 XNOR2_X1 _3031_ (.A(_1717_),
    .B(_1635_),
    .ZN(net72));
 NAND3_X1 _3032_ (.A1(_0153_),
    .A2(_0121_),
    .A3(_0289_),
    .ZN(_0517_));
 NAND2_X1 _3033_ (.A1(net83),
    .A2(_0517_),
    .ZN(_0518_));
 AOI21_X1 _3034_ (.A(_0518_),
    .B1(_0366_),
    .B2(_1687_),
    .ZN(_0519_));
 NAND2_X2 _3035_ (.A1(_0140_),
    .A2(_0281_),
    .ZN(_0520_));
 AOI221_X1 _3036_ (.A(_0520_),
    .B1(_0431_),
    .B2(_0346_),
    .C1(_0405_),
    .C2(_0426_),
    .ZN(_0521_));
 INV_X1 _3037_ (.A(_0521_),
    .ZN(_0522_));
 OAI22_X2 _3038_ (.A1(_0359_),
    .A2(_0413_),
    .B1(_0519_),
    .B2(_0522_),
    .ZN(_0523_));
 OAI211_X2 _3039_ (.A(_0120_),
    .B(_0329_),
    .C1(_0458_),
    .C2(_0461_),
    .ZN(_0524_));
 NOR2_X1 _3040_ (.A1(_1656_),
    .A2(_1660_),
    .ZN(_0525_));
 NOR2_X1 _3041_ (.A1(_1683_),
    .A2(_1671_),
    .ZN(_0526_));
 MUX2_X2 _3042_ (.A(_0525_),
    .B(_0526_),
    .S(_0126_),
    .Z(_0527_));
 OAI21_X1 _3043_ (.A(_0527_),
    .B1(_0451_),
    .B2(_0452_),
    .ZN(_0528_));
 OAI21_X1 _3044_ (.A(_0353_),
    .B1(_0464_),
    .B2(_0465_),
    .ZN(_0529_));
 AND3_X1 _3045_ (.A1(net82),
    .A2(_0126_),
    .A3(_0508_),
    .ZN(_0530_));
 AOI21_X1 _3046_ (.A(_0158_),
    .B1(_0116_),
    .B2(_0068_),
    .ZN(_0531_));
 MUX2_X1 _3047_ (.A(_0531_),
    .B(_0378_),
    .S(_0065_),
    .Z(_0532_));
 OAI21_X1 _3048_ (.A(_0391_),
    .B1(_0530_),
    .B2(_0532_),
    .ZN(_0533_));
 NAND4_X2 _3049_ (.A1(_0524_),
    .A2(_0528_),
    .A3(_0529_),
    .A4(_0533_),
    .ZN(_0534_));
 OAI33_X1 _3050_ (.A1(_0235_),
    .A2(_0454_),
    .A3(_0456_),
    .B1(_0476_),
    .B2(_0478_),
    .B3(_0199_),
    .ZN(_0535_));
 NOR2_X1 _3051_ (.A1(_0481_),
    .A2(_0482_),
    .ZN(_0536_));
 NOR2_X1 _3052_ (.A1(_0473_),
    .A2(_0474_),
    .ZN(_0537_));
 AOI221_X2 _3053_ (.A(_0535_),
    .B1(_0536_),
    .B2(_0353_),
    .C1(_0363_),
    .C2(_0537_),
    .ZN(_0538_));
 MUX2_X1 _3054_ (.A(_0534_),
    .B(_0538_),
    .S(_0153_),
    .Z(_0539_));
 NOR2_X1 _3055_ (.A1(net83),
    .A2(_0539_),
    .ZN(_0540_));
 OAI33_X1 _3056_ (.A1(_0235_),
    .A2(_0469_),
    .A3(_0470_),
    .B1(_0498_),
    .B2(_0499_),
    .B3(_0180_),
    .ZN(_0541_));
 NOR2_X1 _3057_ (.A1(_0494_),
    .A2(_0495_),
    .ZN(_0542_));
 NOR2_X1 _3058_ (.A1(_0491_),
    .A2(_0492_),
    .ZN(_0543_));
 AOI221_X2 _3059_ (.A(_0541_),
    .B1(_0542_),
    .B2(_0363_),
    .C1(_0527_),
    .C2(_0543_),
    .ZN(_0544_));
 AOI21_X1 _3060_ (.A(_1660_),
    .B1(_0081_),
    .B2(_1700_),
    .ZN(_0545_));
 NOR2_X1 _3061_ (.A1(_0126_),
    .A2(_0545_),
    .ZN(_0546_));
 NAND2_X1 _3062_ (.A1(_1700_),
    .A2(_0502_),
    .ZN(_0547_));
 NAND2_X1 _3063_ (.A1(_0192_),
    .A2(_0547_),
    .ZN(_0548_));
 AOI21_X1 _3064_ (.A(_0546_),
    .B1(_0548_),
    .B2(_0126_),
    .ZN(_0549_));
 NOR3_X1 _3065_ (.A1(_0193_),
    .A2(_0487_),
    .A3(_0488_),
    .ZN(_0550_));
 NOR3_X2 _3066_ (.A1(_0120_),
    .A2(_0549_),
    .A3(_0550_),
    .ZN(_0551_));
 MUX2_X1 _3067_ (.A(_0544_),
    .B(_0551_),
    .S(_0153_),
    .Z(_0552_));
 OAI21_X1 _3068_ (.A(_0447_),
    .B1(_0552_),
    .B2(_0151_),
    .ZN(_0553_));
 NOR2_X1 _3069_ (.A1(_0540_),
    .A2(_0553_),
    .ZN(_0554_));
 NOR2_X1 _3070_ (.A1(_0523_),
    .A2(_0554_),
    .ZN(_0555_));
 AND2_X1 _3071_ (.A1(_0523_),
    .A2(_0554_),
    .ZN(_1721_));
 NOR3_X1 _3072_ (.A1(_1701_),
    .A2(_1704_),
    .A3(_0164_),
    .ZN(_0556_));
 NAND3_X1 _3073_ (.A1(_0137_),
    .A2(_0139_),
    .A3(_0556_),
    .ZN(_0557_));
 AND4_X1 _3074_ (.A1(_1693_),
    .A2(_1686_),
    .A3(_0193_),
    .A4(_0357_),
    .ZN(_0558_));
 NOR3_X2 _3075_ (.A1(_0520_),
    .A2(_0557_),
    .A3(_0558_),
    .ZN(_0559_));
 NAND2_X1 _3076_ (.A1(net83),
    .A2(_0559_),
    .ZN(_0560_));
 OAI221_X1 _3077_ (.A(_1573_),
    .B1(_0021_),
    .B2(_0329_),
    .C1(_0357_),
    .C2(_0027_),
    .ZN(_0561_));
 TAPCELL_X1 PHY_12 ();
 OAI21_X1 _3079_ (.A(_0021_),
    .B1(_0329_),
    .B2(_1568_),
    .ZN(_0563_));
 NAND3_X1 _3080_ (.A1(_1558_),
    .A2(_0020_),
    .A3(_0161_),
    .ZN(_0564_));
 NAND3_X1 _3081_ (.A1(_1563_),
    .A2(_0005_),
    .A3(_0357_),
    .ZN(_0565_));
 NAND3_X1 _3082_ (.A1(_0193_),
    .A2(_0564_),
    .A3(_0565_),
    .ZN(_0566_));
 NAND3_X1 _3083_ (.A1(_1563_),
    .A2(_0021_),
    .A3(_0161_),
    .ZN(_0567_));
 NAND3_X1 _3084_ (.A1(_1568_),
    .A2(_0006_),
    .A3(_0357_),
    .ZN(_0568_));
 NAND3_X1 _3085_ (.A1(_0329_),
    .A2(_0567_),
    .A3(_0568_),
    .ZN(_0569_));
 NAND2_X1 _3086_ (.A1(_0566_),
    .A2(_0569_),
    .ZN(_0570_));
 AOI221_X1 _3087_ (.A(_0561_),
    .B1(_0563_),
    .B2(_0357_),
    .C1(_0121_),
    .C2(_0570_),
    .ZN(_0571_));
 MUX2_X1 _3088_ (.A(_1568_),
    .B(_0020_),
    .S(_0357_),
    .Z(_0572_));
 NOR2_X1 _3089_ (.A1(_0329_),
    .A2(_0572_),
    .ZN(_0573_));
 MUX2_X1 _3090_ (.A(_0027_),
    .B(_0030_),
    .S(_0161_),
    .Z(_0574_));
 NAND2_X1 _3091_ (.A1(_1578_),
    .A2(_0574_),
    .ZN(_0575_));
 AOI21_X1 _3092_ (.A(_0573_),
    .B1(_0575_),
    .B2(_0329_),
    .ZN(_0576_));
 AOI221_X1 _3093_ (.A(_0560_),
    .B1(_0571_),
    .B2(_0576_),
    .C1(_1687_),
    .C2(_0121_),
    .ZN(_0577_));
 OAI21_X1 _3094_ (.A(_0527_),
    .B1(_0487_),
    .B2(_0488_),
    .ZN(_0578_));
 OR2_X1 _3095_ (.A1(_0121_),
    .A2(_0503_),
    .ZN(_0579_));
 OAI21_X1 _3096_ (.A(_0391_),
    .B1(_0498_),
    .B2(_0499_),
    .ZN(_0580_));
 AND3_X1 _3097_ (.A1(_0578_),
    .A2(_0579_),
    .A3(_0580_),
    .ZN(_0581_));
 AND4_X1 _3098_ (.A1(_0308_),
    .A2(_0371_),
    .A3(_0412_),
    .A4(_0581_),
    .ZN(_0582_));
 OAI33_X1 _3099_ (.A1(_0199_),
    .A2(_0469_),
    .A3(_0470_),
    .B1(_0481_),
    .B2(_0482_),
    .B3(_0235_),
    .ZN(_0583_));
 AOI221_X2 _3100_ (.A(_0583_),
    .B1(_0542_),
    .B2(_0353_),
    .C1(_0363_),
    .C2(_0543_),
    .ZN(_0584_));
 NAND2_X1 _3101_ (.A1(_0238_),
    .A2(_0404_),
    .ZN(_0585_));
 NOR3_X1 _3102_ (.A1(_0384_),
    .A2(_0584_),
    .A3(_0585_),
    .ZN(_0586_));
 OR2_X1 _3103_ (.A1(_0451_),
    .A2(_0452_),
    .ZN(_0587_));
 OR2_X1 _3104_ (.A1(_0458_),
    .A2(_0461_),
    .ZN(_0588_));
 AOI222_X2 _3105_ (.A1(_0363_),
    .A2(_0587_),
    .B1(_0588_),
    .B2(_0353_),
    .C1(_0512_),
    .C2(_0527_),
    .ZN(_0589_));
 NAND3_X1 _3106_ (.A1(_0405_),
    .A2(_0196_),
    .A3(_0589_),
    .ZN(_0590_));
 NOR2_X1 _3107_ (.A1(_0399_),
    .A2(_0590_),
    .ZN(_0591_));
 NOR3_X1 _3108_ (.A1(_0582_),
    .A2(_0586_),
    .A3(_0591_),
    .ZN(_0592_));
 OAI33_X1 _3109_ (.A1(_0235_),
    .A2(_0464_),
    .A3(_0465_),
    .B1(_0473_),
    .B2(_0474_),
    .B3(_0180_),
    .ZN(_0593_));
 NOR3_X1 _3110_ (.A1(_0199_),
    .A2(_0454_),
    .A3(_0456_),
    .ZN(_0594_));
 NOR4_X1 _3111_ (.A1(_0121_),
    .A2(_0193_),
    .A3(_0476_),
    .A4(_0478_),
    .ZN(_0595_));
 NOR3_X1 _3112_ (.A1(_0593_),
    .A2(_0594_),
    .A3(_0595_),
    .ZN(_0596_));
 NOR3_X1 _3113_ (.A1(_0154_),
    .A2(_0393_),
    .A3(_0596_),
    .ZN(_0597_));
 AOI21_X1 _3114_ (.A(_0520_),
    .B1(_0597_),
    .B2(_0273_),
    .ZN(_0598_));
 AND3_X1 _3115_ (.A1(_1700_),
    .A2(_0125_),
    .A3(_0558_),
    .ZN(_0599_));
 AOI221_X1 _3116_ (.A(_0577_),
    .B1(_0592_),
    .B2(_0598_),
    .C1(_0599_),
    .C2(_0447_),
    .ZN(_0600_));
 TAPCELL_X1 PHY_11 ();
 MUX2_X1 _3118_ (.A(_1558_),
    .B(_1563_),
    .S(_0161_),
    .Z(_0602_));
 NOR2_X1 _3119_ (.A1(_0301_),
    .A2(_0329_),
    .ZN(_0603_));
 MUX2_X1 _3120_ (.A(_1563_),
    .B(_1568_),
    .S(_0161_),
    .Z(_0604_));
 NOR2_X1 _3121_ (.A1(_0017_),
    .A2(_0193_),
    .ZN(_0605_));
 AOI221_X1 _3122_ (.A(_1687_),
    .B1(_0602_),
    .B2(_0603_),
    .C1(_0604_),
    .C2(_0605_),
    .ZN(_0606_));
 MUX2_X1 _3123_ (.A(_0072_),
    .B(_0266_),
    .S(_0161_),
    .Z(_0607_));
 MUX2_X1 _3124_ (.A(_0048_),
    .B(_0049_),
    .S(_0161_),
    .Z(_0608_));
 NAND2_X1 _3125_ (.A1(_1588_),
    .A2(_0608_),
    .ZN(_0609_));
 MUX2_X1 _3126_ (.A(_0575_),
    .B(_0609_),
    .S(_0329_),
    .Z(_0610_));
 NOR4_X1 _3127_ (.A1(_0029_),
    .A2(_0606_),
    .A3(_0607_),
    .A4(_0610_),
    .ZN(_0611_));
 NOR2_X1 _3128_ (.A1(_0001_),
    .A2(_0161_),
    .ZN(_0612_));
 AOI21_X1 _3129_ (.A(_0612_),
    .B1(_0161_),
    .B2(_1553_),
    .ZN(_0613_));
 OR4_X1 _3130_ (.A1(_0284_),
    .A2(_0010_),
    .A3(_0329_),
    .A4(_0613_),
    .ZN(_0614_));
 NAND3_X1 _3131_ (.A1(_1553_),
    .A2(_0006_),
    .A3(_0161_),
    .ZN(_0615_));
 NAND3_X1 _3132_ (.A1(_0005_),
    .A2(_0014_),
    .A3(_0357_),
    .ZN(_0616_));
 AOI21_X1 _3133_ (.A(_0008_),
    .B1(_0615_),
    .B2(_0616_),
    .ZN(_0617_));
 NAND2_X1 _3134_ (.A1(_0329_),
    .A2(_0617_),
    .ZN(_0618_));
 NAND2_X1 _3135_ (.A1(_0005_),
    .A2(_0161_),
    .ZN(_0619_));
 NAND2_X1 _3136_ (.A1(_1553_),
    .A2(_0357_),
    .ZN(_0620_));
 AOI221_X2 _3137_ (.A(_0570_),
    .B1(_0614_),
    .B2(_0618_),
    .C1(_0619_),
    .C2(_0620_),
    .ZN(_0621_));
 NAND2_X1 _3138_ (.A1(_0153_),
    .A2(_0120_),
    .ZN(_0622_));
 MUX2_X1 _3139_ (.A(_0044_),
    .B(_0061_),
    .S(_0357_),
    .Z(_0623_));
 AOI21_X1 _3140_ (.A(_0329_),
    .B1(_0608_),
    .B2(_1588_),
    .ZN(_0624_));
 OAI21_X1 _3141_ (.A(_1598_),
    .B1(_0055_),
    .B2(_0161_),
    .ZN(_0625_));
 AOI21_X1 _3142_ (.A(_0625_),
    .B1(_0161_),
    .B2(_0043_),
    .ZN(_0626_));
 NOR2_X1 _3143_ (.A1(_0193_),
    .A2(_0626_),
    .ZN(_0627_));
 NOR4_X2 _3144_ (.A1(_0088_),
    .A2(_0623_),
    .A3(_0624_),
    .A4(_0627_),
    .ZN(_0628_));
 OAI221_X1 _3145_ (.A(_0611_),
    .B1(_0621_),
    .B2(_0622_),
    .C1(_0628_),
    .C2(_0120_),
    .ZN(_0629_));
 NAND3_X1 _3146_ (.A1(net83),
    .A2(_0559_),
    .A3(_0629_),
    .ZN(_0630_));
 NAND2_X1 _3147_ (.A1(_1603_),
    .A2(_0040_),
    .ZN(_0631_));
 NAND2_X1 _3148_ (.A1(_0329_),
    .A2(_0161_),
    .ZN(_0632_));
 AOI221_X1 _3149_ (.A(_0631_),
    .B1(_0632_),
    .B2(_0043_),
    .C1(_0625_),
    .C2(_0193_),
    .ZN(_0633_));
 OR2_X1 _3150_ (.A1(_0405_),
    .A2(_0633_),
    .ZN(_0634_));
 NAND2_X1 _3151_ (.A1(_0120_),
    .A2(_0283_),
    .ZN(_0635_));
 OAI21_X1 _3152_ (.A(_0035_),
    .B1(_0039_),
    .B2(_0161_),
    .ZN(_0636_));
 AOI221_X2 _3153_ (.A(_1614_),
    .B1(_0193_),
    .B2(_0636_),
    .C1(_0632_),
    .C2(_1611_),
    .ZN(_0637_));
 OAI221_X1 _3154_ (.A(_0634_),
    .B1(_0628_),
    .B2(_0635_),
    .C1(_0637_),
    .C2(_0121_),
    .ZN(_0638_));
 AOI21_X1 _3155_ (.A(_0523_),
    .B1(_0638_),
    .B2(_0559_),
    .ZN(_0639_));
 AND3_X1 _3156_ (.A1(_0600_),
    .A2(_0630_),
    .A3(_0639_),
    .ZN(_0640_));
 NOR3_X1 _3157_ (.A1(_0555_),
    .A2(_1721_),
    .A3(_0640_),
    .ZN(_0641_));
 NOR2_X1 _3158_ (.A1(_0151_),
    .A2(_0310_),
    .ZN(_0642_));
 NAND2_X1 _3159_ (.A1(_0153_),
    .A2(_0148_),
    .ZN(_0643_));
 NAND2_X1 _3160_ (.A1(net84),
    .A2(_0281_),
    .ZN(_0644_));
 OAI22_X2 _3161_ (.A1(_0589_),
    .A2(_0643_),
    .B1(_0644_),
    .B2(_0581_),
    .ZN(_0645_));
 MUX2_X1 _3162_ (.A(_0596_),
    .B(_0584_),
    .S(_0153_),
    .Z(_0646_));
 NOR2_X1 _3163_ (.A1(net83),
    .A2(_0520_),
    .ZN(_0647_));
 AOI22_X4 _3164_ (.A1(_0642_),
    .A2(_0645_),
    .B1(_0646_),
    .B2(_0647_),
    .ZN(_0648_));
 OAI33_X1 _3165_ (.A1(_0235_),
    .A2(_0494_),
    .A3(_0495_),
    .B1(_0498_),
    .B2(_0499_),
    .B3(_0199_),
    .ZN(_0649_));
 NOR4_X1 _3166_ (.A1(_0121_),
    .A2(_0193_),
    .A3(_0487_),
    .A4(_0488_),
    .ZN(_0650_));
 NAND2_X1 _3167_ (.A1(_0177_),
    .A2(_0547_),
    .ZN(_0651_));
 MUX2_X1 _3168_ (.A(_0179_),
    .B(_0651_),
    .S(_0126_),
    .Z(_0652_));
 OAI21_X1 _3169_ (.A(_0652_),
    .B1(_0147_),
    .B2(_0146_),
    .ZN(_0653_));
 OR4_X1 _3170_ (.A1(_0384_),
    .A2(_0649_),
    .A3(_0650_),
    .A4(_0653_),
    .ZN(_0654_));
 OR3_X1 _3171_ (.A1(_0329_),
    .A2(_0451_),
    .A3(_0452_),
    .ZN(_0655_));
 NAND3_X1 _3172_ (.A1(_0329_),
    .A2(_0509_),
    .A3(_0511_),
    .ZN(_0656_));
 NAND4_X1 _3173_ (.A1(_0327_),
    .A2(_0344_),
    .A3(_0655_),
    .A4(_0656_),
    .ZN(_0657_));
 AOI21_X1 _3174_ (.A(_0310_),
    .B1(_0654_),
    .B2(_0657_),
    .ZN(_0658_));
 OAI33_X1 _3175_ (.A1(_0235_),
    .A2(_0473_),
    .A3(_0474_),
    .B1(_0491_),
    .B2(_0492_),
    .B3(_0180_),
    .ZN(_0659_));
 NOR3_X1 _3176_ (.A1(_0199_),
    .A2(_0481_),
    .A3(_0482_),
    .ZN(_0660_));
 NOR4_X1 _3177_ (.A1(_0121_),
    .A2(_0193_),
    .A3(_0469_),
    .A4(_0470_),
    .ZN(_0661_));
 OR3_X2 _3178_ (.A1(_0659_),
    .A2(_0660_),
    .A3(_0661_),
    .ZN(_0662_));
 NOR4_X1 _3179_ (.A1(_0121_),
    .A2(_0193_),
    .A3(_0454_),
    .A4(_0456_),
    .ZN(_0663_));
 NOR3_X1 _3180_ (.A1(_0180_),
    .A2(_0476_),
    .A3(_0478_),
    .ZN(_0664_));
 NOR3_X1 _3181_ (.A1(_0235_),
    .A2(_0458_),
    .A3(_0461_),
    .ZN(_0665_));
 NOR3_X1 _3182_ (.A1(_0199_),
    .A2(_0464_),
    .A3(_0465_),
    .ZN(_0666_));
 OR4_X2 _3183_ (.A1(_0663_),
    .A2(_0664_),
    .A3(_0665_),
    .A4(_0666_),
    .ZN(_0667_));
 OAI22_X2 _3184_ (.A1(_0408_),
    .A2(_0662_),
    .B1(_0667_),
    .B2(_0406_),
    .ZN(_0668_));
 OAI21_X2 _3185_ (.A(_1723_),
    .B1(_0658_),
    .B2(_0668_),
    .ZN(_0669_));
 NOR4_X4 _3186_ (.A1(_0444_),
    .A2(_0449_),
    .A3(_0648_),
    .A4(_0669_),
    .ZN(_1733_));
 AOI21_X1 _3187_ (.A(_0281_),
    .B1(_0534_),
    .B2(_0153_),
    .ZN(_0670_));
 NOR2_X1 _3188_ (.A1(net83),
    .A2(_0281_),
    .ZN(_0671_));
 AOI221_X1 _3189_ (.A(_0151_),
    .B1(_0279_),
    .B2(_0280_),
    .C1(_0551_),
    .C2(net85),
    .ZN(_0672_));
 OAI221_X1 _3190_ (.A(_0140_),
    .B1(_0154_),
    .B2(_0544_),
    .C1(_0538_),
    .C2(_0283_),
    .ZN(_0673_));
 OR4_X2 _3191_ (.A1(_0670_),
    .A2(_0671_),
    .A3(_0672_),
    .A4(_0673_),
    .ZN(_0674_));
 AOI211_X2 _3192_ (.A(_0436_),
    .B(_0674_),
    .C1(_0281_),
    .C2(_0440_),
    .ZN(_0675_));
 OAI221_X2 _3193_ (.A(_0148_),
    .B1(_0427_),
    .B2(_0467_),
    .C1(_0513_),
    .C2(_0384_),
    .ZN(_0676_));
 AOI21_X1 _3194_ (.A(_0148_),
    .B1(_0420_),
    .B2(_0504_),
    .ZN(_0677_));
 OAI221_X2 _3195_ (.A(_0677_),
    .B1(_0501_),
    .B2(_0154_),
    .C1(_0283_),
    .C2(_0484_),
    .ZN(_0678_));
 NAND3_X2 _3196_ (.A1(_0140_),
    .A2(_0676_),
    .A3(_0678_),
    .ZN(_0679_));
 NOR3_X2 _3197_ (.A1(_0430_),
    .A2(_0434_),
    .A3(_0679_),
    .ZN(_0680_));
 INV_X1 _3198_ (.A(_0652_),
    .ZN(_0681_));
 OR3_X1 _3199_ (.A1(_0681_),
    .A2(_0649_),
    .A3(_0650_),
    .ZN(_0682_));
 NOR2_X1 _3200_ (.A1(_0408_),
    .A2(_0682_),
    .ZN(_0683_));
 NAND2_X1 _3201_ (.A1(_0655_),
    .A2(_0656_),
    .ZN(_0684_));
 OAI21_X1 _3202_ (.A(_1687_),
    .B1(_0121_),
    .B2(_0684_),
    .ZN(_0685_));
 NAND2_X2 _3203_ (.A1(_1693_),
    .A2(_0148_),
    .ZN(_0686_));
 NOR3_X1 _3204_ (.A1(_0310_),
    .A2(_0686_),
    .A3(_0667_),
    .ZN(_0687_));
 AOI21_X1 _3205_ (.A(_0683_),
    .B1(_0685_),
    .B2(_0687_),
    .ZN(_0688_));
 NAND2_X1 _3206_ (.A1(_0281_),
    .A2(_0405_),
    .ZN(_0689_));
 NOR2_X1 _3207_ (.A1(_0689_),
    .A2(_0662_),
    .ZN(_0690_));
 NOR2_X1 _3208_ (.A1(_0421_),
    .A2(_0684_),
    .ZN(_0691_));
 OAI21_X1 _3209_ (.A(_0140_),
    .B1(_0690_),
    .B2(_0691_),
    .ZN(_0692_));
 AOI21_X2 _3210_ (.A(_0425_),
    .B1(_0688_),
    .B2(_0692_),
    .ZN(_0693_));
 NAND4_X4 _3211_ (.A1(_1733_),
    .A2(_0675_),
    .A3(_0680_),
    .A4(_0693_),
    .ZN(_0694_));
 NOR2_X1 _3212_ (.A1(_0689_),
    .A2(_0581_),
    .ZN(_0695_));
 OAI21_X1 _3213_ (.A(_0151_),
    .B1(net84),
    .B2(_0589_),
    .ZN(_0696_));
 AOI21_X1 _3214_ (.A(_0695_),
    .B1(_0696_),
    .B2(_0148_),
    .ZN(_0697_));
 OAI21_X1 _3215_ (.A(_0140_),
    .B1(_0646_),
    .B2(_0151_),
    .ZN(_0698_));
 NOR2_X1 _3216_ (.A1(_0697_),
    .A2(_0698_),
    .ZN(_0699_));
 NAND2_X1 _3217_ (.A1(_1760_),
    .A2(_0699_),
    .ZN(_0700_));
 NOR3_X1 _3218_ (.A1(_0310_),
    .A2(_0148_),
    .A3(_0283_),
    .ZN(_0701_));
 AND2_X1 _3219_ (.A1(_0701_),
    .A2(_0584_),
    .ZN(_0702_));
 NOR2_X1 _3220_ (.A1(_0408_),
    .A2(_0581_),
    .ZN(_0703_));
 OR3_X1 _3221_ (.A1(_0593_),
    .A2(_0594_),
    .A3(_0595_),
    .ZN(_0704_));
 OAI22_X1 _3222_ (.A1(_0413_),
    .A2(_0704_),
    .B1(_0589_),
    .B2(_0415_),
    .ZN(_0705_));
 OAI33_X1 _3223_ (.A1(_0414_),
    .A2(_0416_),
    .A3(_0417_),
    .B1(_0702_),
    .B2(_0703_),
    .B3(_0705_),
    .ZN(_0706_));
 OAI21_X1 _3224_ (.A(_0671_),
    .B1(_0684_),
    .B2(_0622_),
    .ZN(_0707_));
 OAI21_X1 _3225_ (.A(_0281_),
    .B1(_0283_),
    .B2(_0682_),
    .ZN(_0708_));
 NAND3_X1 _3226_ (.A1(_0140_),
    .A2(_0707_),
    .A3(_0708_),
    .ZN(_0709_));
 MUX2_X1 _3227_ (.A(_0662_),
    .B(_0667_),
    .S(net84),
    .Z(_0710_));
 AND2_X1 _3228_ (.A1(net83),
    .A2(_0710_),
    .ZN(_0711_));
 NOR3_X1 _3229_ (.A1(_0706_),
    .A2(_0709_),
    .A3(_0711_),
    .ZN(_0712_));
 NOR2_X1 _3230_ (.A1(_0310_),
    .A2(_0407_),
    .ZN(_0713_));
 AOI22_X1 _3231_ (.A1(_0701_),
    .A2(_0544_),
    .B1(_0551_),
    .B2(_0713_),
    .ZN(_0714_));
 AOI22_X1 _3232_ (.A1(_0395_),
    .A2(_0534_),
    .B1(_0538_),
    .B2(_0394_),
    .ZN(_0715_));
 NAND2_X1 _3233_ (.A1(_0714_),
    .A2(_0715_),
    .ZN(_0716_));
 AND2_X1 _3234_ (.A1(_1749_),
    .A2(_0716_),
    .ZN(_0717_));
 MUX2_X1 _3235_ (.A(_0505_),
    .B(_0513_),
    .S(_0148_),
    .Z(_0718_));
 OAI222_X2 _3236_ (.A1(_0686_),
    .A2(_0485_),
    .B1(_0501_),
    .B2(_0689_),
    .C1(_0718_),
    .C2(_0154_),
    .ZN(_0719_));
 AND2_X1 _3237_ (.A1(_1752_),
    .A2(_0719_),
    .ZN(_0720_));
 NAND3_X1 _3238_ (.A1(_0712_),
    .A2(_0717_),
    .A3(_0720_),
    .ZN(_0721_));
 NAND2_X1 _3239_ (.A1(_0151_),
    .A2(_0140_),
    .ZN(_0722_));
 AOI21_X1 _3240_ (.A(_0148_),
    .B1(_0551_),
    .B2(net85),
    .ZN(_0723_));
 AND2_X1 _3241_ (.A1(_0153_),
    .A2(_0544_),
    .ZN(_0724_));
 AOI21_X1 _3242_ (.A(_0724_),
    .B1(_0538_),
    .B2(net84),
    .ZN(_0725_));
 OAI33_X1 _3243_ (.A1(_0722_),
    .A2(_0670_),
    .A3(_0723_),
    .B1(_0725_),
    .B2(_0310_),
    .B3(_0686_),
    .ZN(_0726_));
 NOR2_X1 _3244_ (.A1(_0310_),
    .A2(_0686_),
    .ZN(_0727_));
 INV_X1 _3245_ (.A(_0727_),
    .ZN(_0728_));
 NAND2_X1 _3246_ (.A1(_0153_),
    .A2(_0399_),
    .ZN(_0729_));
 MUX2_X1 _3247_ (.A(_0437_),
    .B(_0729_),
    .S(_0148_),
    .Z(_0730_));
 OAI22_X2 _3248_ (.A1(_0728_),
    .A2(_0439_),
    .B1(_0722_),
    .B2(_0730_),
    .ZN(_1764_));
 NAND2_X1 _3249_ (.A1(_0726_),
    .A2(_1764_),
    .ZN(_0731_));
 NAND3_X1 _3250_ (.A1(_0117_),
    .A2(_0140_),
    .A3(_0325_),
    .ZN(_0732_));
 NAND3_X1 _3251_ (.A1(_0151_),
    .A2(_0144_),
    .A3(_0331_),
    .ZN(_0733_));
 OAI21_X1 _3252_ (.A(_0733_),
    .B1(_0144_),
    .B2(_0151_),
    .ZN(_0734_));
 NOR2_X1 _3253_ (.A1(_0151_),
    .A2(_0343_),
    .ZN(_0735_));
 OR4_X1 _3254_ (.A1(_0731_),
    .A2(_0732_),
    .A3(_0734_),
    .A4(_0735_),
    .ZN(_0736_));
 NOR4_X2 _3255_ (.A1(_0694_),
    .A2(_0700_),
    .A3(_0721_),
    .A4(_0736_),
    .ZN(_0737_));
 TAPCELL_X1 PHY_10 ();
 MUX2_X1 _3257_ (.A(_0641_),
    .B(_1724_),
    .S(net81),
    .Z(net49));
 MUX2_X1 _3258_ (.A(_1724_),
    .B(_1727_),
    .S(net81),
    .Z(net60));
 OR2_X1 _3259_ (.A1(_0658_),
    .A2(_0668_),
    .ZN(_0739_));
 XOR2_X1 _3260_ (.A(_1726_),
    .B(_0739_),
    .Z(_0740_));
 MUX2_X1 _3261_ (.A(_1727_),
    .B(_0740_),
    .S(net81),
    .Z(net71));
 MUX2_X1 _3262_ (.A(_0740_),
    .B(_1731_),
    .S(net81),
    .Z(net74));
 XNOR2_X1 _3263_ (.A(_1730_),
    .B(_0648_),
    .ZN(_0741_));
 MUX2_X1 _3264_ (.A(_1731_),
    .B(_0741_),
    .S(net81),
    .Z(net75));
 MUX2_X1 _3265_ (.A(_0741_),
    .B(_1735_),
    .S(net81),
    .Z(net76));
 XNOR2_X1 _3266_ (.A(_1734_),
    .B(_0674_),
    .ZN(_0742_));
 MUX2_X1 _3267_ (.A(_1735_),
    .B(_0742_),
    .S(net81),
    .Z(net77));
 MUX2_X1 _3268_ (.A(_0742_),
    .B(_1739_),
    .S(net81),
    .Z(net78));
 XNOR2_X1 _3269_ (.A(_1738_),
    .B(_0679_),
    .ZN(_0743_));
 MUX2_X1 _3270_ (.A(_1739_),
    .B(_0743_),
    .S(net81),
    .Z(net79));
 AND2_X1 _3271_ (.A1(_1733_),
    .A2(_0675_),
    .ZN(_1736_));
 AND2_X1 _3272_ (.A1(_1736_),
    .A2(_0680_),
    .ZN(_1741_));
 MUX2_X1 _3273_ (.A(_0743_),
    .B(_1743_),
    .S(net81),
    .Z(net80));
 NAND2_X1 _3274_ (.A1(_0688_),
    .A2(_0692_),
    .ZN(_0744_));
 XOR2_X1 _3275_ (.A(_1742_),
    .B(_0744_),
    .Z(_0745_));
 TAPCELL_X1 PHY_9 ();
 MUX2_X1 _3277_ (.A(_1743_),
    .B(_0745_),
    .S(net81),
    .Z(net50));
 MUX2_X1 _3278_ (.A(_0745_),
    .B(_1747_),
    .S(net81),
    .Z(net51));
 OR3_X1 _3279_ (.A1(_0702_),
    .A2(_0703_),
    .A3(_0705_),
    .ZN(_0747_));
 XOR2_X1 _3280_ (.A(_1746_),
    .B(_0747_),
    .Z(_0748_));
 MUX2_X1 _3281_ (.A(_1747_),
    .B(_0748_),
    .S(net81),
    .Z(net52));
 NOR2_X1 _3282_ (.A1(_0694_),
    .A2(_0706_),
    .ZN(_1748_));
 MUX2_X1 _3283_ (.A(_0748_),
    .B(_1751_),
    .S(net81),
    .Z(net53));
 XOR2_X1 _3284_ (.A(_1750_),
    .B(_0716_),
    .Z(_0749_));
 MUX2_X1 _3285_ (.A(_1751_),
    .B(_0749_),
    .S(net81),
    .Z(net54));
 MUX2_X1 _3286_ (.A(_0749_),
    .B(_1755_),
    .S(net81),
    .Z(net55));
 NAND2_X1 _3287_ (.A1(_0140_),
    .A2(_0719_),
    .ZN(_0750_));
 XNOR2_X1 _3288_ (.A(_1754_),
    .B(_0750_),
    .ZN(_0751_));
 MUX2_X1 _3289_ (.A(_1755_),
    .B(_0751_),
    .S(net81),
    .Z(net56));
 AND2_X1 _3290_ (.A1(_0717_),
    .A2(_1748_),
    .ZN(_1753_));
 AND2_X1 _3291_ (.A1(_0720_),
    .A2(_1753_),
    .ZN(_1757_));
 MUX2_X1 _3292_ (.A(_0751_),
    .B(_1759_),
    .S(net81),
    .Z(net57));
 NOR2_X1 _3293_ (.A1(_0709_),
    .A2(_0711_),
    .ZN(_0752_));
 XOR2_X1 _3294_ (.A(_1758_),
    .B(_0752_),
    .Z(_0753_));
 MUX2_X1 _3295_ (.A(_1759_),
    .B(_0753_),
    .S(net81),
    .Z(net58));
 MUX2_X1 _3296_ (.A(_0753_),
    .B(_1763_),
    .S(net81),
    .Z(net59));
 XOR2_X1 _3297_ (.A(_1762_),
    .B(_0699_),
    .Z(_0754_));
 MUX2_X1 _3298_ (.A(_1763_),
    .B(_0754_),
    .S(_0737_),
    .Z(net61));
 NAND3_X1 _3299_ (.A1(_0712_),
    .A2(_0717_),
    .A3(_0720_),
    .ZN(_0755_));
 NOR4_X1 _3300_ (.A1(_0310_),
    .A2(_0345_),
    .A3(_0694_),
    .A4(_0755_),
    .ZN(_1761_));
 AND3_X1 _3301_ (.A1(_1760_),
    .A2(_0699_),
    .A3(_1761_),
    .ZN(_1765_));
 MUX2_X1 _3302_ (.A(_0754_),
    .B(_1767_),
    .S(_0737_),
    .Z(net62));
 XOR2_X1 _3303_ (.A(_1766_),
    .B(_0726_),
    .Z(_0756_));
 MUX2_X1 _3304_ (.A(_1767_),
    .B(_0756_),
    .S(_0737_),
    .Z(net63));
 INV_X1 _3305_ (.A(_1661_),
    .ZN(_1682_));
 NAND2_X1 _3306_ (.A1(net32),
    .A2(net92),
    .ZN(_0757_));
 OAI21_X4 _3307_ (.A(_0757_),
    .B1(net92),
    .B2(_1843_),
    .ZN(_1616_));
 NAND4_X1 _3308_ (.A1(_1657_),
    .A2(_1650_),
    .A3(_1642_),
    .A4(_0068_),
    .ZN(_0758_));
 OR4_X1 _3309_ (.A1(_0111_),
    .A2(_1682_),
    .A3(_1616_),
    .A4(_0758_),
    .ZN(_0759_));
 NOR2_X1 _3310_ (.A1(_1548_),
    .A2(_0759_),
    .ZN(_1615_));
 INV_X1 _3311_ (.A(_1647_),
    .ZN(_1630_));
 INV_X1 _3312_ (.A(_1623_),
    .ZN(net65));
 INV_X1 _3313_ (.A(_1627_),
    .ZN(net66));
 INV_X1 _3314_ (.A(_1636_),
    .ZN(net70));
 NOR2_X1 _3315_ (.A1(_0110_),
    .A2(_0759_),
    .ZN(_1679_));
 XNOR2_X1 _3316_ (.A(_1670_),
    .B(_1646_),
    .ZN(_0760_));
 MUX2_X1 _3317_ (.A(_1645_),
    .B(_0760_),
    .S(_0126_),
    .Z(_1684_));
 INV_X1 _3318_ (.A(_1718_),
    .ZN(_1715_));
 NOR2_X1 _3319_ (.A1(_0449_),
    .A2(_0669_),
    .ZN(_1728_));
 INV_X1 _3320_ (.A(_0694_),
    .ZN(_1744_));
 NOR2_X1 _3321_ (.A1(net92),
    .A2(_1813_),
    .ZN(_0761_));
 TAPCELL_X1 PHY_8 ();
 AOI21_X1 _3323_ (.A(_0761_),
    .B1(net92),
    .B2(net31),
    .ZN(_0763_));
 XNOR2_X1 _3324_ (.A(_1222_),
    .B(_0763_),
    .ZN(_1845_));
 MUX2_X1 _3325_ (.A(net30),
    .B(_1275_),
    .S(_1131_),
    .Z(_0764_));
 XOR2_X2 _3326_ (.A(_1222_),
    .B(_0764_),
    .Z(_1550_));
 MUX2_X1 _3327_ (.A(_1326_),
    .B(_1819_),
    .S(_1131_),
    .Z(_0765_));
 XNOR2_X1 _3328_ (.A(_1222_),
    .B(_0765_),
    .ZN(_1851_));
 NAND2_X1 _3329_ (.A1(net27),
    .A2(net92),
    .ZN(_0766_));
 OAI21_X1 _3330_ (.A(_0766_),
    .B1(_1822_),
    .B2(net92),
    .ZN(_0767_));
 XOR2_X2 _3331_ (.A(_1222_),
    .B(_0767_),
    .Z(_1555_));
 NAND2_X1 _3332_ (.A1(_1196_),
    .A2(_1217_),
    .ZN(_0768_));
 OAI21_X1 _3333_ (.A(_0768_),
    .B1(_1313_),
    .B2(_1196_),
    .ZN(_0769_));
 NAND3_X1 _3334_ (.A1(_1135_),
    .A2(_1184_),
    .A3(_0769_),
    .ZN(_0770_));
 NOR2_X1 _3335_ (.A1(_1139_),
    .A2(_0770_),
    .ZN(_0771_));
 OR2_X1 _3336_ (.A1(net97),
    .A2(_1309_),
    .ZN(_0772_));
 OAI21_X1 _3337_ (.A(_0772_),
    .B1(_1327_),
    .B2(_1196_),
    .ZN(_0773_));
 AND3_X1 _3338_ (.A1(_1317_),
    .A2(_1319_),
    .A3(_1322_),
    .ZN(_0774_));
 MUX2_X1 _3339_ (.A(_0774_),
    .B(_1335_),
    .S(net96),
    .Z(_0775_));
 MUX2_X1 _3340_ (.A(_0773_),
    .B(_0775_),
    .S(_1135_),
    .Z(_0776_));
 AOI21_X2 _3341_ (.A(_0771_),
    .B1(_0776_),
    .B2(_1402_),
    .ZN(_0777_));
 NOR2_X1 _3342_ (.A1(_1191_),
    .A2(_0777_),
    .ZN(_0778_));
 XNOR2_X1 _3343_ (.A(_1202_),
    .B(_0778_),
    .ZN(_1857_));
 NAND2_X1 _3344_ (.A1(_1209_),
    .A2(_1385_),
    .ZN(_0779_));
 XNOR2_X2 _3345_ (.A(_1379_),
    .B(_0779_),
    .ZN(_1560_));
 MUX2_X1 _3346_ (.A(net24),
    .B(_1303_),
    .S(_1131_),
    .Z(_0780_));
 XOR2_X1 _3347_ (.A(_1222_),
    .B(_0780_),
    .Z(_1863_));
 MUX2_X1 _3348_ (.A(net23),
    .B(_1304_),
    .S(_1131_),
    .Z(_0781_));
 XOR2_X2 _3349_ (.A(_1222_),
    .B(_0781_),
    .Z(_1565_));
 NAND2_X1 _3350_ (.A1(net22),
    .A2(net90),
    .ZN(_0782_));
 OAI21_X1 _3351_ (.A(_0782_),
    .B1(_1837_),
    .B2(net90),
    .ZN(_0783_));
 XOR2_X1 _3352_ (.A(_1222_),
    .B(_0783_),
    .Z(_1869_));
 AND2_X1 _3353_ (.A1(_1196_),
    .A2(_1340_),
    .ZN(_0784_));
 NAND2_X1 _3354_ (.A1(net93),
    .A2(net20),
    .ZN(_0785_));
 NOR2_X1 _3355_ (.A1(net90),
    .A2(_0785_),
    .ZN(_0786_));
 OAI21_X1 _3356_ (.A(_1184_),
    .B1(_0784_),
    .B2(_0786_),
    .ZN(_0787_));
 NOR2_X1 _3357_ (.A1(_1134_),
    .A2(_0787_),
    .ZN(_0788_));
 AND2_X1 _3358_ (.A1(_1342_),
    .A2(_1343_),
    .ZN(_0789_));
 NAND2_X1 _3359_ (.A1(net96),
    .A2(_0789_),
    .ZN(_0790_));
 NAND2_X1 _3360_ (.A1(_1346_),
    .A2(_1347_),
    .ZN(_0791_));
 OAI21_X1 _3361_ (.A(_0790_),
    .B1(_0791_),
    .B2(net96),
    .ZN(_0792_));
 NOR2_X1 _3362_ (.A1(_1135_),
    .A2(_1355_),
    .ZN(_0793_));
 AOI21_X1 _3363_ (.A(_0788_),
    .B1(_0792_),
    .B2(_0793_),
    .ZN(_0794_));
 AOI21_X1 _3364_ (.A(_1138_),
    .B1(_1187_),
    .B2(_0794_),
    .ZN(_0795_));
 NAND2_X1 _3365_ (.A1(_0769_),
    .A2(_0793_),
    .ZN(_0796_));
 NAND2_X1 _3366_ (.A1(_1196_),
    .A2(_1309_),
    .ZN(_0797_));
 NOR2_X1 _3367_ (.A1(net29),
    .A2(net90),
    .ZN(_0798_));
 AOI21_X1 _3368_ (.A(_0798_),
    .B1(_1819_),
    .B2(net90),
    .ZN(_0799_));
 OAI211_X2 _3369_ (.A(_1135_),
    .B(_0797_),
    .C1(_0799_),
    .C2(_1196_),
    .ZN(_0800_));
 OAI21_X1 _3370_ (.A(_0796_),
    .B1(_0800_),
    .B2(_1355_),
    .ZN(_0801_));
 OAI21_X1 _3371_ (.A(_0795_),
    .B1(_0801_),
    .B2(_1187_),
    .ZN(_0802_));
 OAI21_X1 _3372_ (.A(_1196_),
    .B1(net25),
    .B2(net90),
    .ZN(_0803_));
 AND2_X1 _3373_ (.A1(_1301_),
    .A2(_1330_),
    .ZN(_0804_));
 OAI22_X1 _3374_ (.A1(_1196_),
    .A2(_1350_),
    .B1(_0803_),
    .B2(_0804_),
    .ZN(_0805_));
 MUX2_X1 _3375_ (.A(_0775_),
    .B(_0805_),
    .S(_1135_),
    .Z(_0806_));
 AND2_X1 _3376_ (.A1(_1184_),
    .A2(_0806_),
    .ZN(_0807_));
 NAND3_X1 _3377_ (.A1(_1138_),
    .A2(_1187_),
    .A3(_0807_),
    .ZN(_0808_));
 AOI21_X1 _3378_ (.A(_1208_),
    .B1(_0802_),
    .B2(_0808_),
    .ZN(_0809_));
 XNOR2_X1 _3379_ (.A(_1202_),
    .B(_0809_),
    .ZN(_1877_));
 NAND2_X1 _3380_ (.A1(net19),
    .A2(net91),
    .ZN(_0810_));
 XNOR2_X2 _3381_ (.A(_1222_),
    .B(_0810_),
    .ZN(_1575_));
 NAND2_X1 _3382_ (.A1(net18),
    .A2(net91),
    .ZN(_0811_));
 XNOR2_X1 _3383_ (.A(_1222_),
    .B(_0811_),
    .ZN(_1883_));
 NAND2_X1 _3384_ (.A1(net47),
    .A2(net91),
    .ZN(_0812_));
 XNOR2_X1 _3385_ (.A(_1222_),
    .B(_0812_),
    .ZN(_1891_));
 AND2_X1 _3386_ (.A1(_1409_),
    .A2(_1414_),
    .ZN(_1895_));
 NAND3_X1 _3387_ (.A1(_1135_),
    .A2(_1402_),
    .A3(_0769_),
    .ZN(_0813_));
 MUX2_X1 _3388_ (.A(net48),
    .B(net47),
    .S(net97),
    .Z(_0814_));
 MUX2_X1 _3389_ (.A(net46),
    .B(net45),
    .S(net97),
    .Z(_0815_));
 MUX2_X1 _3390_ (.A(_0814_),
    .B(_0815_),
    .S(_1135_),
    .Z(_0816_));
 NAND2_X1 _3391_ (.A1(_1365_),
    .A2(_0816_),
    .ZN(_0817_));
 NOR2_X1 _3392_ (.A1(_1138_),
    .A2(_0817_),
    .ZN(_0818_));
 NAND2_X1 _3393_ (.A1(_1196_),
    .A2(net19),
    .ZN(_0819_));
 INV_X1 _3394_ (.A(net18),
    .ZN(_0820_));
 OAI21_X1 _3395_ (.A(_0819_),
    .B1(_0820_),
    .B2(_1196_),
    .ZN(_0821_));
 NAND3_X1 _3396_ (.A1(_1135_),
    .A2(_1365_),
    .A3(_0821_),
    .ZN(_0822_));
 OAI21_X1 _3397_ (.A(_0822_),
    .B1(_0787_),
    .B2(_1135_),
    .ZN(_0823_));
 AOI21_X1 _3398_ (.A(_0818_),
    .B1(_0823_),
    .B2(_1138_),
    .ZN(_0824_));
 OAI22_X1 _3399_ (.A1(_1417_),
    .A2(_0813_),
    .B1(_0824_),
    .B2(_1191_),
    .ZN(_0825_));
 OR2_X1 _3400_ (.A1(_1134_),
    .A2(_0775_),
    .ZN(_0826_));
 OAI21_X1 _3401_ (.A(_0826_),
    .B1(_0773_),
    .B2(_1135_),
    .ZN(_0827_));
 OAI21_X1 _3402_ (.A(_1138_),
    .B1(_1355_),
    .B2(_0827_),
    .ZN(_0828_));
 MUX2_X1 _3403_ (.A(_0792_),
    .B(_0805_),
    .S(_1134_),
    .Z(_0829_));
 AOI21_X1 _3404_ (.A(_1138_),
    .B1(_1184_),
    .B2(_0829_),
    .ZN(_0830_));
 NOR2_X1 _3405_ (.A1(_1307_),
    .A2(_0830_),
    .ZN(_0831_));
 AOI21_X1 _3406_ (.A(_0825_),
    .B1(_0828_),
    .B2(_0831_),
    .ZN(_0832_));
 XNOR2_X1 _3407_ (.A(_1379_),
    .B(_0832_),
    .ZN(_1899_));
 NAND2_X1 _3408_ (.A1(net43),
    .A2(net91),
    .ZN(_0833_));
 XNOR2_X1 _3409_ (.A(_1222_),
    .B(_0833_),
    .ZN(_1907_));
 NOR2_X1 _3410_ (.A1(_1196_),
    .A2(_1456_),
    .ZN(_0834_));
 MUX2_X1 _3411_ (.A(net44),
    .B(net42),
    .S(_1135_),
    .Z(_0835_));
 AOI21_X1 _3412_ (.A(_0834_),
    .B1(_0835_),
    .B2(_1196_),
    .ZN(_0836_));
 OAI22_X1 _3413_ (.A1(_1139_),
    .A2(_0817_),
    .B1(_0836_),
    .B2(_1461_),
    .ZN(_0837_));
 NAND2_X1 _3414_ (.A1(_1209_),
    .A2(_0837_),
    .ZN(_0838_));
 INV_X1 _3415_ (.A(_0823_),
    .ZN(_0839_));
 NAND2_X1 _3416_ (.A1(_1184_),
    .A2(_0829_),
    .ZN(_0840_));
 MUX2_X1 _3417_ (.A(_0839_),
    .B(_0840_),
    .S(_1138_),
    .Z(_0841_));
 OAI221_X2 _3418_ (.A(_0838_),
    .B1(_0777_),
    .B2(_1417_),
    .C1(_1307_),
    .C2(_0841_),
    .ZN(_0842_));
 XNOR2_X1 _3419_ (.A(_1202_),
    .B(_0842_),
    .ZN(_1915_));
 NOR2_X1 _3420_ (.A1(_1135_),
    .A2(_0815_),
    .ZN(_0843_));
 AND2_X1 _3421_ (.A1(_1196_),
    .A2(net44),
    .ZN(_0844_));
 AOI21_X1 _3422_ (.A(_0844_),
    .B1(net43),
    .B2(net95),
    .ZN(_0845_));
 AOI21_X1 _3423_ (.A(_0843_),
    .B1(_0845_),
    .B2(_1135_),
    .ZN(_0846_));
 NAND2_X1 _3424_ (.A1(_1365_),
    .A2(_0846_),
    .ZN(_0847_));
 TAPCELL_X1 PHY_7 ();
 MUX2_X1 _3426_ (.A(net39),
    .B(net17),
    .S(_1135_),
    .Z(_0849_));
 AND2_X1 _3427_ (.A1(net94),
    .A2(_0849_),
    .ZN(_0850_));
 AOI21_X1 _3428_ (.A(_0850_),
    .B1(_1459_),
    .B2(_1196_),
    .ZN(_0851_));
 OAI22_X1 _3429_ (.A1(_1139_),
    .A2(_0847_),
    .B1(_0851_),
    .B2(_1461_),
    .ZN(_0852_));
 NOR3_X1 _3430_ (.A1(_1134_),
    .A2(_1384_),
    .A3(_1417_),
    .ZN(_0853_));
 AOI22_X1 _3431_ (.A1(_1209_),
    .A2(_0852_),
    .B1(_0853_),
    .B2(_0773_),
    .ZN(_0854_));
 MUX2_X1 _3432_ (.A(_0821_),
    .B(_0814_),
    .S(_1135_),
    .Z(_0855_));
 NAND2_X1 _3433_ (.A1(_1365_),
    .A2(_0855_),
    .ZN(_0856_));
 MUX2_X1 _3434_ (.A(_0794_),
    .B(_0856_),
    .S(_1139_),
    .Z(_0857_));
 OAI21_X1 _3435_ (.A(_0854_),
    .B1(_0857_),
    .B2(_1307_),
    .ZN(_0858_));
 AOI21_X1 _3436_ (.A(_1417_),
    .B1(_0796_),
    .B2(_1138_),
    .ZN(_0859_));
 NAND2_X1 _3437_ (.A1(_1184_),
    .A2(_0806_),
    .ZN(_0860_));
 NAND2_X1 _3438_ (.A1(_1139_),
    .A2(_0860_),
    .ZN(_0861_));
 AOI21_X1 _3439_ (.A(_0858_),
    .B1(_0859_),
    .B2(_0861_),
    .ZN(_0862_));
 XNOR2_X1 _3440_ (.A(_1379_),
    .B(_0862_),
    .ZN(_1923_));
 NAND2_X1 _3441_ (.A1(_1365_),
    .A2(_1446_),
    .ZN(_0863_));
 AND2_X1 _3442_ (.A1(net95),
    .A2(net28),
    .ZN(_0864_));
 AOI22_X1 _3443_ (.A1(_1196_),
    .A2(_0849_),
    .B1(_0864_),
    .B2(_1134_),
    .ZN(_0865_));
 OAI22_X1 _3444_ (.A1(_1139_),
    .A2(_0863_),
    .B1(_1461_),
    .B2(_0865_),
    .ZN(_0866_));
 NOR3_X2 _3445_ (.A1(_1142_),
    .A2(_1187_),
    .A3(_1189_),
    .ZN(_0867_));
 AOI22_X1 _3446_ (.A1(_1209_),
    .A2(_0866_),
    .B1(_0867_),
    .B2(_1219_),
    .ZN(_0868_));
 NOR2_X1 _3447_ (.A1(_1355_),
    .A2(_1417_),
    .ZN(_0869_));
 INV_X1 _3448_ (.A(_0869_),
    .ZN(_0870_));
 MUX2_X1 _3449_ (.A(_1436_),
    .B(_1407_),
    .S(_1138_),
    .Z(_0871_));
 OAI221_X2 _3450_ (.A(_0868_),
    .B1(_0870_),
    .B2(_0871_),
    .C1(_1399_),
    .C2(_1307_),
    .ZN(_0872_));
 XNOR2_X2 _3451_ (.A(_1202_),
    .B(_0872_),
    .ZN(_1605_));
 AND2_X1 _3452_ (.A1(_1196_),
    .A2(net28),
    .ZN(_0873_));
 AOI21_X1 _3453_ (.A(_0873_),
    .B1(net17),
    .B2(net94),
    .ZN(_0874_));
 OAI22_X1 _3454_ (.A1(_1139_),
    .A2(_0836_),
    .B1(_0874_),
    .B2(_1429_),
    .ZN(_0875_));
 NAND3_X1 _3455_ (.A1(_1209_),
    .A2(_1365_),
    .A3(_0875_),
    .ZN(_0876_));
 NAND2_X1 _3456_ (.A1(_1139_),
    .A2(_1453_),
    .ZN(_0877_));
 OAI221_X2 _3457_ (.A(_0876_),
    .B1(_0840_),
    .B2(_0877_),
    .C1(_1307_),
    .C2(_0824_),
    .ZN(_0878_));
 INV_X1 _3458_ (.A(_0813_),
    .ZN(_0879_));
 NOR2_X1 _3459_ (.A1(_1384_),
    .A2(_1417_),
    .ZN(_0880_));
 AOI221_X2 _3460_ (.A(_0878_),
    .B1(_0867_),
    .B2(_0879_),
    .C1(_0776_),
    .C2(_0880_),
    .ZN(_0881_));
 XNOR2_X1 _3461_ (.A(_1379_),
    .B(_0881_),
    .ZN(_1610_));
 AOI21_X1 _3462_ (.A(_1189_),
    .B1(_1946_),
    .B2(_1947_),
    .ZN(_1929_));
 NAND3_X1 _3463_ (.A1(_1937_),
    .A2(_1139_),
    .A3(_0867_),
    .ZN(_0882_));
 NAND3_X1 _3464_ (.A1(_1184_),
    .A2(_1929_),
    .A3(_0882_),
    .ZN(_0883_));
 XNOR2_X1 _3465_ (.A(_1948_),
    .B(_1189_),
    .ZN(_0884_));
 XNOR2_X1 _3466_ (.A(_1770_),
    .B(_1931_),
    .ZN(_0885_));
 XNOR2_X1 _3467_ (.A(_1537_),
    .B(_0885_),
    .ZN(_0886_));
 OR3_X2 _3468_ (.A1(_1932_),
    .A2(net91),
    .A3(_0886_),
    .ZN(_0887_));
 TAPCELL_X1 PHY_6 ();
 TAPCELL_X1 PHY_5 ();
 TAPCELL_X1 PHY_4 ();
 TAPCELL_X1 PHY_3 ();
 INV_X1 _3473_ (.A(net42),
    .ZN(_0892_));
 OAI21_X1 _3474_ (.A(_1444_),
    .B1(_0892_),
    .B2(net94),
    .ZN(_0893_));
 AOI21_X1 _3475_ (.A(_0893_),
    .B1(net44),
    .B2(net94),
    .ZN(_0894_));
 NOR3_X1 _3476_ (.A1(net39),
    .A2(_1936_),
    .A3(_0873_),
    .ZN(_0895_));
 AOI221_X1 _3477_ (.A(_1945_),
    .B1(_1936_),
    .B2(_0894_),
    .C1(_0895_),
    .C2(_1442_),
    .ZN(_0896_));
 INV_X1 _3478_ (.A(_0896_),
    .ZN(_0897_));
 TAPCELL_X1 PHY_2 ();
 NAND2_X1 _3480_ (.A1(_1945_),
    .A2(_1936_),
    .ZN(_0899_));
 NOR2_X1 _3481_ (.A1(net17),
    .A2(_0864_),
    .ZN(_0900_));
 OAI21_X1 _3482_ (.A(_0897_),
    .B1(_0899_),
    .B2(_0900_),
    .ZN(_0901_));
 INV_X2 _3483_ (.A(net89),
    .ZN(_0902_));
 TAPCELL_X1 PHY_1 ();
 AND2_X1 _3485_ (.A1(net95),
    .A2(net46),
    .ZN(_0904_));
 NOR4_X1 _3486_ (.A1(net45),
    .A2(_0902_),
    .A3(_0904_),
    .A4(_0844_),
    .ZN(_0905_));
 AOI21_X1 _3487_ (.A(_0905_),
    .B1(_0894_),
    .B2(_0902_),
    .ZN(_0906_));
 NOR3_X1 _3488_ (.A1(net93),
    .A2(net19),
    .A3(net47),
    .ZN(_0907_));
 NOR2_X1 _3489_ (.A1(net20),
    .A2(net48),
    .ZN(_0908_));
 AOI21_X1 _3490_ (.A(_0907_),
    .B1(_0908_),
    .B2(net93),
    .ZN(_0909_));
 NOR3_X1 _3491_ (.A1(net93),
    .A2(net48),
    .A3(net45),
    .ZN(_0910_));
 NOR2_X1 _3492_ (.A1(net18),
    .A2(net46),
    .ZN(_0911_));
 AOI21_X1 _3493_ (.A(_0910_),
    .B1(_0911_),
    .B2(net93),
    .ZN(_0912_));
 MUX2_X1 _3494_ (.A(_0909_),
    .B(_0912_),
    .S(_0902_),
    .Z(_0913_));
 INV_X1 _3495_ (.A(net48),
    .ZN(_0914_));
 OR2_X1 _3496_ (.A1(net47),
    .A2(net89),
    .ZN(_0915_));
 AOI21_X1 _3497_ (.A(_0915_),
    .B1(net46),
    .B2(_1196_),
    .ZN(_0916_));
 NAND2_X1 _3498_ (.A1(_0914_),
    .A2(_0916_),
    .ZN(_0917_));
 NAND2_X1 _3499_ (.A1(net95),
    .A2(net89),
    .ZN(_0918_));
 OR2_X1 _3500_ (.A1(net19),
    .A2(net18),
    .ZN(_0919_));
 NOR3_X1 _3501_ (.A1(net18),
    .A2(net48),
    .A3(_0902_),
    .ZN(_0920_));
 NOR2_X1 _3502_ (.A1(_0916_),
    .A2(_0920_),
    .ZN(_0921_));
 OAI221_X2 _3503_ (.A(_0917_),
    .B1(_0918_),
    .B2(_0919_),
    .C1(net93),
    .C2(_0921_),
    .ZN(_0922_));
 NOR3_X1 _3504_ (.A1(net93),
    .A2(net46),
    .A3(net43),
    .ZN(_0923_));
 NOR2_X1 _3505_ (.A1(net48),
    .A2(net44),
    .ZN(_0924_));
 AOI21_X1 _3506_ (.A(_0923_),
    .B1(_0924_),
    .B2(net93),
    .ZN(_0925_));
 NOR3_X1 _3507_ (.A1(net47),
    .A2(_0902_),
    .A3(_0925_),
    .ZN(_0926_));
 NOR3_X1 _3508_ (.A1(net93),
    .A2(net44),
    .A3(net39),
    .ZN(_0927_));
 NOR2_X1 _3509_ (.A1(net46),
    .A2(net42),
    .ZN(_0928_));
 AOI21_X1 _3510_ (.A(_0927_),
    .B1(_0928_),
    .B2(net93),
    .ZN(_0929_));
 NOR3_X1 _3511_ (.A1(net45),
    .A2(_1936_),
    .A3(_0929_),
    .ZN(_0930_));
 NOR2_X1 _3512_ (.A1(net17),
    .A2(_1936_),
    .ZN(_0931_));
 NOR2_X1 _3513_ (.A1(net39),
    .A2(net28),
    .ZN(_0932_));
 AOI21_X1 _3514_ (.A(_0931_),
    .B1(_0932_),
    .B2(_1936_),
    .ZN(_0933_));
 NOR2_X1 _3515_ (.A1(net95),
    .A2(_0933_),
    .ZN(_0934_));
 OAI33_X1 _3516_ (.A1(net28),
    .A2(net17),
    .A3(net89),
    .B1(_0918_),
    .B2(net42),
    .B3(net39),
    .ZN(_0935_));
 OAI221_X1 _3517_ (.A(_0922_),
    .B1(_0926_),
    .B2(_0930_),
    .C1(_0934_),
    .C2(_0935_),
    .ZN(_0936_));
 MUX2_X1 _3518_ (.A(_0913_),
    .B(_0936_),
    .S(_1945_),
    .Z(_0937_));
 NOR3_X1 _3519_ (.A1(_0901_),
    .A2(_0906_),
    .A3(_0937_),
    .ZN(_0938_));
 OAI21_X1 _3520_ (.A(_1949_),
    .B1(_0887_),
    .B2(_0938_),
    .ZN(_0939_));
 MUX2_X1 _3521_ (.A(net18),
    .B(net19),
    .S(net93),
    .Z(_0940_));
 NAND2_X1 _3522_ (.A1(_0902_),
    .A2(_0940_),
    .ZN(_0941_));
 AOI21_X1 _3523_ (.A(_0887_),
    .B1(_0922_),
    .B2(_0941_),
    .ZN(_0942_));
 AOI21_X1 _3524_ (.A(net28),
    .B1(_1936_),
    .B2(net42),
    .ZN(_0943_));
 NOR2_X1 _3525_ (.A1(_1196_),
    .A2(_0943_),
    .ZN(_0944_));
 NOR2_X1 _3526_ (.A1(_0902_),
    .A2(_0932_),
    .ZN(_0945_));
 NOR3_X1 _3527_ (.A1(net17),
    .A2(_0944_),
    .A3(_0945_),
    .ZN(_0946_));
 NOR3_X1 _3528_ (.A1(net88),
    .A2(_0887_),
    .A3(_0946_),
    .ZN(_0947_));
 XNOR2_X2 _3529_ (.A(_1944_),
    .B(_1205_),
    .ZN(_0948_));
 AOI21_X1 _3530_ (.A(_0942_),
    .B1(_0947_),
    .B2(_0948_),
    .ZN(_0949_));
 NOR2_X1 _3531_ (.A1(net88),
    .A2(_0949_),
    .ZN(_0950_));
 NOR2_X1 _3532_ (.A1(_0939_),
    .A2(_0950_),
    .ZN(_0951_));
 XNOR2_X1 _3533_ (.A(_1182_),
    .B(_0885_),
    .ZN(_0952_));
 NOR2_X1 _3534_ (.A1(_1932_),
    .A2(_0952_),
    .ZN(_0953_));
 NAND2_X1 _3535_ (.A1(net89),
    .A2(_0953_),
    .ZN(_0954_));
 INV_X1 _3536_ (.A(net20),
    .ZN(_0955_));
 OAI21_X1 _3537_ (.A(_1196_),
    .B1(_0955_),
    .B2(net90),
    .ZN(_0956_));
 OAI21_X1 _3538_ (.A(_0956_),
    .B1(_1340_),
    .B2(_1196_),
    .ZN(_0957_));
 OR2_X1 _3539_ (.A1(_0954_),
    .A2(_0957_),
    .ZN(_0958_));
 NOR2_X1 _3540_ (.A1(_1196_),
    .A2(_0902_),
    .ZN(_0959_));
 NAND4_X1 _3541_ (.A1(_1346_),
    .A2(_1347_),
    .A3(_0959_),
    .A4(_0953_),
    .ZN(_0960_));
 OR2_X1 _3542_ (.A1(_1932_),
    .A2(_0952_),
    .ZN(_0961_));
 AOI221_X1 _3543_ (.A(_0902_),
    .B1(_1342_),
    .B2(_1343_),
    .C1(_1340_),
    .C2(_1196_),
    .ZN(_0962_));
 NAND2_X1 _3544_ (.A1(_0955_),
    .A2(_0819_),
    .ZN(_0963_));
 AOI221_X1 _3545_ (.A(net89),
    .B1(_1131_),
    .B2(_0963_),
    .C1(_1340_),
    .C2(net96),
    .ZN(_0964_));
 OR3_X1 _3546_ (.A1(_0961_),
    .A2(_0962_),
    .A3(_0964_),
    .ZN(_0965_));
 AND3_X1 _3547_ (.A1(_0958_),
    .A2(_0960_),
    .A3(_0965_),
    .ZN(_0966_));
 OAI21_X1 _3548_ (.A(_0951_),
    .B1(_0966_),
    .B2(net88),
    .ZN(_0967_));
 INV_X1 _3549_ (.A(_0887_),
    .ZN(_0968_));
 MUX2_X1 _3550_ (.A(net44),
    .B(net46),
    .S(_1936_),
    .Z(_0969_));
 MUX2_X1 _3551_ (.A(net45),
    .B(net47),
    .S(_1936_),
    .Z(_0970_));
 MUX2_X1 _3552_ (.A(_0969_),
    .B(_0970_),
    .S(net94),
    .Z(_0971_));
 MUX2_X1 _3553_ (.A(net28),
    .B(net42),
    .S(_1936_),
    .Z(_0972_));
 MUX2_X1 _3554_ (.A(net39),
    .B(net43),
    .S(_1936_),
    .Z(_0973_));
 MUX2_X1 _3555_ (.A(_0972_),
    .B(_0973_),
    .S(net94),
    .Z(_0974_));
 MUX2_X1 _3556_ (.A(_0971_),
    .B(_0974_),
    .S(_1945_),
    .Z(_0975_));
 AND3_X1 _3557_ (.A1(_1949_),
    .A2(_0968_),
    .A3(_0975_),
    .ZN(_0976_));
 OR3_X1 _3558_ (.A1(_0948_),
    .A2(_0947_),
    .A3(_0976_),
    .ZN(_0977_));
 NOR2_X1 _3559_ (.A1(_0935_),
    .A2(_0934_),
    .ZN(_0978_));
 MUX2_X1 _3560_ (.A(_0906_),
    .B(_0978_),
    .S(_1945_),
    .Z(_0979_));
 NOR2_X1 _3561_ (.A1(_0901_),
    .A2(_0979_),
    .ZN(_0980_));
 NOR2_X1 _3562_ (.A1(_0887_),
    .A2(_0980_),
    .ZN(_0981_));
 OAI21_X1 _3563_ (.A(_0948_),
    .B1(_0947_),
    .B2(_0981_),
    .ZN(_0982_));
 INV_X1 _3564_ (.A(_0982_),
    .ZN(_0983_));
 OAI221_X1 _3565_ (.A(_0884_),
    .B1(_0967_),
    .B2(_0977_),
    .C1(_0983_),
    .C2(_1949_),
    .ZN(_0984_));
 OAI21_X1 _3566_ (.A(_1202_),
    .B1(_0883_),
    .B2(_0984_),
    .ZN(_0985_));
 OR3_X1 _3567_ (.A1(_0774_),
    .A2(_1331_),
    .A3(_1335_),
    .ZN(_0986_));
 AND2_X1 _3568_ (.A1(_1309_),
    .A2(_1313_),
    .ZN(_0987_));
 NOR3_X1 _3569_ (.A1(net20),
    .A2(net47),
    .A3(net17),
    .ZN(_0988_));
 NOR4_X1 _3570_ (.A1(net46),
    .A2(net44),
    .A3(net43),
    .A4(net42),
    .ZN(_0989_));
 NOR3_X1 _3571_ (.A1(net48),
    .A2(net45),
    .A3(_0919_),
    .ZN(_0990_));
 NAND4_X1 _3572_ (.A1(_0988_),
    .A2(_0989_),
    .A3(_0932_),
    .A4(_0990_),
    .ZN(_0991_));
 AND2_X1 _3573_ (.A1(_1131_),
    .A2(_0991_),
    .ZN(_0992_));
 NOR4_X1 _3574_ (.A1(_1217_),
    .A2(_1340_),
    .A3(_0789_),
    .A4(_0992_),
    .ZN(_0993_));
 AND3_X1 _3575_ (.A1(_0791_),
    .A2(_1350_),
    .A3(_0993_),
    .ZN(_0994_));
 NAND3_X1 _3576_ (.A1(_1327_),
    .A2(_0987_),
    .A3(_0994_),
    .ZN(_0995_));
 OAI21_X1 _3577_ (.A(_0883_),
    .B1(_0986_),
    .B2(_0995_),
    .ZN(_0996_));
 MUX2_X1 _3578_ (.A(_1202_),
    .B(_0985_),
    .S(_0996_),
    .Z(_0997_));
 OR3_X1 _3579_ (.A1(_1202_),
    .A2(_0883_),
    .A3(_0984_),
    .ZN(_0998_));
 OR2_X1 _3580_ (.A1(_1379_),
    .A2(_0883_),
    .ZN(_0999_));
 NOR2_X1 _3581_ (.A1(net88),
    .A2(_0953_),
    .ZN(_1000_));
 AOI21_X1 _3582_ (.A(_1196_),
    .B1(net89),
    .B2(_1217_),
    .ZN(_1001_));
 AOI22_X1 _3583_ (.A1(_1196_),
    .A2(_1323_),
    .B1(_1309_),
    .B2(_1001_),
    .ZN(_1002_));
 NOR3_X1 _3584_ (.A1(net88),
    .A2(_0799_),
    .A3(_1002_),
    .ZN(_1003_));
 AOI211_X2 _3585_ (.A(_1324_),
    .B(_1335_),
    .C1(_1331_),
    .C2(_1196_),
    .ZN(_1004_));
 MUX2_X1 _3586_ (.A(_0987_),
    .B(_1004_),
    .S(_0902_),
    .Z(_1005_));
 NAND3_X1 _3587_ (.A1(_0958_),
    .A2(_0960_),
    .A3(_0965_),
    .ZN(_1006_));
 NOR2_X1 _3588_ (.A1(net89),
    .A2(_0784_),
    .ZN(_1007_));
 AOI21_X1 _3589_ (.A(_0961_),
    .B1(_1007_),
    .B2(_0790_),
    .ZN(_1008_));
 NOR2_X1 _3590_ (.A1(net96),
    .A2(_0902_),
    .ZN(_1009_));
 AOI22_X1 _3591_ (.A1(_1350_),
    .A2(_0959_),
    .B1(_1009_),
    .B2(_0791_),
    .ZN(_1010_));
 INV_X1 _3592_ (.A(_0941_),
    .ZN(_1011_));
 AOI221_X1 _3593_ (.A(_1006_),
    .B1(_1008_),
    .B2(_1010_),
    .C1(_1011_),
    .C2(_0968_),
    .ZN(_1012_));
 AOI221_X1 _3594_ (.A(_1000_),
    .B1(_1003_),
    .B2(_1005_),
    .C1(net88),
    .C2(_1012_),
    .ZN(_1013_));
 INV_X1 _3595_ (.A(net17),
    .ZN(_1014_));
 NOR4_X1 _3596_ (.A1(_1014_),
    .A2(net88),
    .A3(_0887_),
    .A4(_0918_),
    .ZN(_1015_));
 AOI21_X1 _3597_ (.A(_1949_),
    .B1(_0948_),
    .B2(_1015_),
    .ZN(_1016_));
 NAND3_X1 _3598_ (.A1(net89),
    .A2(_0785_),
    .A3(_0819_),
    .ZN(_1017_));
 AOI21_X1 _3599_ (.A(net89),
    .B1(net18),
    .B2(net93),
    .ZN(_1018_));
 OAI21_X1 _3600_ (.A(_1018_),
    .B1(_0914_),
    .B2(net93),
    .ZN(_1019_));
 NAND4_X1 _3601_ (.A1(net88),
    .A2(_0968_),
    .A3(_1017_),
    .A4(_1019_),
    .ZN(_1020_));
 NAND2_X1 _3602_ (.A1(_1008_),
    .A2(_1010_),
    .ZN(_1021_));
 AOI21_X1 _3603_ (.A(_1016_),
    .B1(_1020_),
    .B2(_1021_),
    .ZN(_1022_));
 NAND2_X1 _3604_ (.A1(_0968_),
    .A2(_0975_),
    .ZN(_1023_));
 AND2_X1 _3605_ (.A1(_0948_),
    .A2(_1023_),
    .ZN(_1024_));
 NAND4_X1 _3606_ (.A1(_0791_),
    .A2(_1350_),
    .A3(_1344_),
    .A4(_0948_),
    .ZN(_1025_));
 OAI21_X1 _3607_ (.A(net89),
    .B1(_1350_),
    .B2(net96),
    .ZN(_1026_));
 AOI22_X1 _3608_ (.A1(net96),
    .A2(_1331_),
    .B1(_1025_),
    .B2(_1026_),
    .ZN(_1027_));
 OAI221_X1 _3609_ (.A(_1024_),
    .B1(_1027_),
    .B2(_0961_),
    .C1(_0954_),
    .C2(_1004_),
    .ZN(_1028_));
 NOR4_X1 _3610_ (.A1(_0967_),
    .A2(_1013_),
    .A3(_1022_),
    .A4(_1028_),
    .ZN(_1029_));
 MUX2_X1 _3611_ (.A(_0998_),
    .B(_0999_),
    .S(_1029_),
    .Z(_1030_));
 AND2_X1 _3612_ (.A1(_0997_),
    .A2(_1030_),
    .ZN(_1612_));
 INV_X1 _3613_ (.A(_1507_),
    .ZN(_1554_));
 OR2_X1 _3614_ (.A1(_1865_),
    .A2(_1506_),
    .ZN(_1559_));
 INV_X1 _3615_ (.A(_1872_),
    .ZN(_1031_));
 OAI21_X1 _3616_ (.A(_1504_),
    .B1(_1503_),
    .B2(_1031_),
    .ZN(_1564_));
 INV_X1 _3617_ (.A(_1885_),
    .ZN(_1032_));
 AND3_X1 _3618_ (.A1(_1890_),
    .A2(_1482_),
    .A3(_1485_),
    .ZN(_1033_));
 OAI21_X1 _3619_ (.A(_1886_),
    .B1(_1889_),
    .B2(_1033_),
    .ZN(_1034_));
 NAND2_X1 _3620_ (.A1(_1032_),
    .A2(_1034_),
    .ZN(_1574_));
 AND3_X1 _3621_ (.A1(_0726_),
    .A2(_1764_),
    .A3(_1765_),
    .ZN(_1617_));
 INV_X1 _3622_ (.A(_1664_),
    .ZN(_1625_));
 INV_X1 _3623_ (.A(_1713_),
    .ZN(_1035_));
 INV_X1 _3624_ (.A(_1711_),
    .ZN(_1036_));
 NOR2_X1 _3625_ (.A1(_1036_),
    .A2(_1629_),
    .ZN(_1037_));
 OAI21_X1 _3626_ (.A(_1714_),
    .B1(_1710_),
    .B2(_1037_),
    .ZN(_1038_));
 NAND2_X1 _3627_ (.A1(_1035_),
    .A2(_1038_),
    .ZN(_1634_));
 INV_X1 _3628_ (.A(_1519_),
    .ZN(_1523_));
 INV_X1 _3629_ (.A(_1511_),
    .ZN(_1515_));
 INV_X1 _3630_ (.A(_1843_),
    .ZN(_1841_));
 NOR2_X1 _3631_ (.A1(_1191_),
    .A2(_0813_),
    .ZN(_1039_));
 XNOR2_X1 _3632_ (.A(_1202_),
    .B(_1039_),
    .ZN(_1846_));
 NOR3_X1 _3633_ (.A1(_1185_),
    .A2(_1191_),
    .A3(_1315_),
    .ZN(_1040_));
 XNOR2_X2 _3634_ (.A(_1202_),
    .B(_1040_),
    .ZN(_1551_));
 NAND3_X1 _3635_ (.A1(_1139_),
    .A2(_1209_),
    .A3(_0801_),
    .ZN(_1041_));
 XNOR2_X1 _3636_ (.A(_1379_),
    .B(_1041_),
    .ZN(_1852_));
 NOR2_X1 _3637_ (.A1(_1191_),
    .A2(_1435_),
    .ZN(_1042_));
 XNOR2_X2 _3638_ (.A(_1202_),
    .B(_1042_),
    .ZN(_1556_));
 MUX2_X1 _3639_ (.A(_1334_),
    .B(_1825_),
    .S(_1131_),
    .Z(_1043_));
 XNOR2_X1 _3640_ (.A(_1222_),
    .B(_1043_),
    .ZN(_1858_));
 NAND2_X1 _3641_ (.A1(net25),
    .A2(net90),
    .ZN(_1044_));
 OAI21_X1 _3642_ (.A(_1044_),
    .B1(_1828_),
    .B2(net90),
    .ZN(_1045_));
 XOR2_X2 _3643_ (.A(_1222_),
    .B(_1045_),
    .Z(_1561_));
 MUX2_X1 _3644_ (.A(_0801_),
    .B(_0807_),
    .S(_1139_),
    .Z(_1046_));
 NAND2_X1 _3645_ (.A1(_1209_),
    .A2(_1046_),
    .ZN(_1047_));
 XNOR2_X1 _3646_ (.A(_1379_),
    .B(_1047_),
    .ZN(_1864_));
 NOR2_X1 _3647_ (.A1(_1384_),
    .A2(_1407_),
    .ZN(_1048_));
 NAND2_X1 _3648_ (.A1(_1187_),
    .A2(_1404_),
    .ZN(_1049_));
 OAI221_X2 _3649_ (.A(_1190_),
    .B1(_1048_),
    .B2(_1049_),
    .C1(_1219_),
    .C2(_1187_),
    .ZN(_1050_));
 XNOR2_X2 _3650_ (.A(_1379_),
    .B(_1050_),
    .ZN(_1566_));
 AOI21_X1 _3651_ (.A(_1139_),
    .B1(_1184_),
    .B2(_0776_),
    .ZN(_1051_));
 OAI33_X1 _3652_ (.A1(_1138_),
    .A2(_1307_),
    .A3(_0770_),
    .B1(_1051_),
    .B2(_0830_),
    .B3(_1191_),
    .ZN(_1052_));
 XNOR2_X1 _3653_ (.A(_1202_),
    .B(_1052_),
    .ZN(_1870_));
 XNOR2_X1 _3654_ (.A(_1379_),
    .B(_1359_),
    .ZN(_1874_));
 NAND2_X1 _3655_ (.A1(net20),
    .A2(net91),
    .ZN(_1053_));
 XNOR2_X1 _3656_ (.A(_1222_),
    .B(_1053_),
    .ZN(_1878_));
 NOR3_X1 _3657_ (.A1(_1205_),
    .A2(_1437_),
    .A3(_1439_),
    .ZN(_1054_));
 AOI211_X2 _3658_ (.A(_1208_),
    .B(_1054_),
    .C1(_1435_),
    .C2(_1205_),
    .ZN(_1055_));
 XNOR2_X2 _3659_ (.A(_1202_),
    .B(_1055_),
    .ZN(_1576_));
 OAI22_X1 _3660_ (.A1(_1307_),
    .A2(_0777_),
    .B1(_0841_),
    .B2(_1191_),
    .ZN(_1056_));
 XNOR2_X1 _3661_ (.A(_1202_),
    .B(_1056_),
    .ZN(_1884_));
 OR2_X1 _3662_ (.A1(_1205_),
    .A2(_1377_),
    .ZN(_1057_));
 MUX2_X1 _3663_ (.A(_1202_),
    .B(_1362_),
    .S(_1385_),
    .Z(_1058_));
 OAI221_X2 _3664_ (.A(_1057_),
    .B1(_1202_),
    .B2(_1190_),
    .C1(_1187_),
    .C2(_1058_),
    .ZN(_1888_));
 NAND2_X1 _3665_ (.A1(_1187_),
    .A2(_0857_),
    .ZN(_1059_));
 OAI211_X2 _3666_ (.A(_1190_),
    .B(_1059_),
    .C1(_1046_),
    .C2(_1187_),
    .ZN(_1060_));
 XNOR2_X1 _3667_ (.A(_1379_),
    .B(_1060_),
    .ZN(_1892_));
 NAND2_X1 _3668_ (.A1(net45),
    .A2(net91),
    .ZN(_1061_));
 XNOR2_X1 _3669_ (.A(_1222_),
    .B(_1061_),
    .ZN(_1900_));
 XNOR2_X1 _3670_ (.A(_1202_),
    .B(_1427_),
    .ZN(_1904_));
 NOR3_X1 _3671_ (.A1(_1139_),
    .A2(_1191_),
    .A3(_0856_),
    .ZN(_1062_));
 OAI222_X2 _3672_ (.A1(_1417_),
    .A2(_0796_),
    .B1(_0870_),
    .B2(_0800_),
    .C1(_0847_),
    .C2(_1191_),
    .ZN(_1063_));
 INV_X1 _3673_ (.A(_1307_),
    .ZN(_1064_));
 OR2_X1 _3674_ (.A1(_1138_),
    .A2(_0794_),
    .ZN(_1065_));
 OAI21_X1 _3675_ (.A(_1065_),
    .B1(_0860_),
    .B2(_1139_),
    .ZN(_1066_));
 AOI221_X2 _3676_ (.A(_1062_),
    .B1(_1063_),
    .B2(_1139_),
    .C1(_1064_),
    .C2(_1066_),
    .ZN(_1067_));
 XNOR2_X1 _3677_ (.A(_1379_),
    .B(_1067_),
    .ZN(_1908_));
 XNOR2_X1 _3678_ (.A(_1202_),
    .B(_1450_),
    .ZN(_1912_));
 NAND2_X1 _3679_ (.A1(net39),
    .A2(net91),
    .ZN(_1068_));
 XNOR2_X1 _3680_ (.A(_1222_),
    .B(_1068_),
    .ZN(_1916_));
 XNOR2_X1 _3681_ (.A(_1379_),
    .B(_1463_),
    .ZN(_1920_));
 NAND2_X1 _3682_ (.A1(net17),
    .A2(net91),
    .ZN(_1069_));
 XNOR2_X1 _3683_ (.A(_1222_),
    .B(_1069_),
    .ZN(_1924_));
 FA_X1 _3684_ (.A(net33),
    .B(_1510_),
    .CI(_1511_),
    .CO(_1512_),
    .S(_1513_));
 FA_X1 _3685_ (.A(_1514_),
    .B(_1515_),
    .CI(_1516_),
    .CO(_1517_),
    .S(_1518_));
 FA_X1 _3686_ (.A(net34),
    .B(_1519_),
    .CI(_1512_),
    .CO(_1520_),
    .S(_1521_));
 FA_X1 _3687_ (.A(_1522_),
    .B(_1523_),
    .CI(_1517_),
    .CO(_1524_),
    .S(_1525_));
 FA_X1 _3688_ (.A(_1526_),
    .B(_1527_),
    .CI(_1528_),
    .CO(_1529_),
    .S(_1530_));
 FA_X1 _3689_ (.A(net36),
    .B(_1531_),
    .CI(_1532_),
    .CO(_1533_),
    .S(_1534_));
 FA_X1 _3690_ (.A(net38),
    .B(_1535_),
    .CI(_1536_),
    .CO(_1537_),
    .S(_1538_));
 FA_X1 _3691_ (.A(_1539_),
    .B(_1540_),
    .CI(_1541_),
    .CO(_1542_),
    .S(_1543_));
 FA_X1 _3692_ (.A(_1544_),
    .B(_1545_),
    .CI(_1546_),
    .CO(_1547_),
    .S(_1548_));
 FA_X1 _3693_ (.A(_1549_),
    .B(_1550_),
    .CI(_1551_),
    .CO(_1552_),
    .S(_1553_));
 FA_X1 _3694_ (.A(_1554_),
    .B(_1555_),
    .CI(_1556_),
    .CO(_1557_),
    .S(_1558_));
 FA_X1 _3695_ (.A(_1559_),
    .B(_1560_),
    .CI(_1561_),
    .CO(_1562_),
    .S(_1563_));
 FA_X1 _3696_ (.A(_1564_),
    .B(_1565_),
    .CI(_1566_),
    .CO(_1567_),
    .S(_1568_));
 FA_X1 _3697_ (.A(_1569_),
    .B(_1570_),
    .CI(_1571_),
    .CO(_1572_),
    .S(_1573_));
 FA_X1 _3698_ (.A(_1574_),
    .B(_1575_),
    .CI(_1576_),
    .CO(_1577_),
    .S(_1578_));
 FA_X1 _3699_ (.A(_1579_),
    .B(_1580_),
    .CI(_1581_),
    .CO(_1582_),
    .S(_1583_));
 FA_X1 _3700_ (.A(_1584_),
    .B(_1585_),
    .CI(_1586_),
    .CO(_1587_),
    .S(_1588_));
 FA_X1 _3701_ (.A(_1589_),
    .B(_1590_),
    .CI(_1591_),
    .CO(_1592_),
    .S(_1593_));
 FA_X1 _3702_ (.A(_1594_),
    .B(_1595_),
    .CI(_1596_),
    .CO(_1597_),
    .S(_1598_));
 FA_X1 _3703_ (.A(_1599_),
    .B(_1600_),
    .CI(_1601_),
    .CO(_1602_),
    .S(_1603_));
 FA_X1 _3704_ (.A(_1604_),
    .B(_1605_),
    .CI(_1222_),
    .CO(_1607_),
    .S(_1608_));
 FA_X1 _3705_ (.A(_1609_),
    .B(_1610_),
    .CI(_1222_),
    .CO(_1604_),
    .S(_1611_));
 FA_X1 _3706_ (.A(_1612_),
    .B(_1222_),
    .CI(_1613_),
    .CO(_1609_),
    .S(_1614_));
 FA_X1 _3707_ (.A(_1615_),
    .B(_1616_),
    .CI(_1617_),
    .CO(_1618_),
    .S(_1619_));
 FA_X1 _3708_ (.A(_1620_),
    .B(_1621_),
    .CI(_1618_),
    .CO(_1622_),
    .S(_1623_));
 FA_X1 _3709_ (.A(_1624_),
    .B(_1625_),
    .CI(_1622_),
    .CO(_1626_),
    .S(_1627_));
 FA_X1 _3710_ (.A(_1628_),
    .B(_1629_),
    .CI(_1630_),
    .CO(_1631_),
    .S(net68));
 FA_X1 _3711_ (.A(_1632_),
    .B(_1633_),
    .CI(_1634_),
    .CO(_1635_),
    .S(_1636_));
 HA_X1 _3712_ (.A(_1637_),
    .B(_1638_),
    .CO(_1639_),
    .S(_1640_));
 HA_X1 _3713_ (.A(_1641_),
    .B(_1642_),
    .CO(_1643_),
    .S(_1644_));
 HA_X1 _3714_ (.A(_1645_),
    .B(_1646_),
    .CO(_1647_),
    .S(_1648_));
 HA_X1 _3715_ (.A(_1649_),
    .B(_1650_),
    .CO(_1651_),
    .S(_1652_));
 HA_X1 _3716_ (.A(_1653_),
    .B(_1654_),
    .CO(_1655_),
    .S(_1624_));
 HA_X1 _3717_ (.A(_1656_),
    .B(_1657_),
    .CO(_1658_),
    .S(_1659_));
 HA_X1 _3718_ (.A(_1660_),
    .B(_1661_),
    .CO(_1662_),
    .S(_1663_));
 HA_X1 _3719_ (.A(_1660_),
    .B(_1661_),
    .CO(_1664_),
    .S(_1665_));
 HA_X1 _3720_ (.A(_1616_),
    .B(_0065_),
    .CO(_1667_),
    .S(_1668_));
 HA_X1 _3721_ (.A(_1669_),
    .B(_1654_),
    .CO(_1670_),
    .S(_1671_));
 HA_X1 _3722_ (.A(_1672_),
    .B(_1673_),
    .CO(_1674_),
    .S(_1675_));
 HA_X1 _3723_ (.A(_1676_),
    .B(_1638_),
    .CO(_1677_),
    .S(_1678_));
 HA_X1 _3724_ (.A(_1679_),
    .B(_1616_),
    .CO(_1680_),
    .S(_1681_));
 HA_X1 _3725_ (.A(_1680_),
    .B(_1682_),
    .CO(_1669_),
    .S(_1683_));
 HA_X1 _3726_ (.A(_1684_),
    .B(_0120_),
    .CO(_1686_),
    .S(_1687_));
 HA_X1 _3727_ (.A(_1684_),
    .B(_0121_),
    .CO(_1689_),
    .S(_1690_));
 HA_X1 _3728_ (.A(_1689_),
    .B(_1691_),
    .CO(_1692_),
    .S(_1693_));
 HA_X1 _3729_ (.A(_1694_),
    .B(_1695_),
    .CO(_1696_),
    .S(_1697_));
 HA_X1 _3730_ (.A(_1698_),
    .B(_1699_),
    .CO(_1700_),
    .S(_1701_));
 HA_X1 _3731_ (.A(_1702_),
    .B(_1703_),
    .CO(_1704_),
    .S(_1705_));
 HA_X1 _3732_ (.A(_0065_),
    .B(_1619_),
    .CO(_1621_),
    .S(net64));
 HA_X1 _3733_ (.A(_1624_),
    .B(_1625_),
    .CO(_1706_),
    .S(_1707_));
 HA_X1 _3734_ (.A(_1648_),
    .B(_1655_),
    .CO(_1708_),
    .S(_1709_));
 HA_X1 _3735_ (.A(_1640_),
    .B(_1647_),
    .CO(_1710_),
    .S(_1711_));
 HA_X1 _3736_ (.A(_0068_),
    .B(_1639_),
    .CO(_1713_),
    .S(_1714_));
 HA_X1 _3737_ (.A(_1715_),
    .B(_1632_),
    .CO(_1716_),
    .S(_1717_));
 HA_X1 _3738_ (.A(_1718_),
    .B(_1673_),
    .CO(_1719_),
    .S(_1720_));
 HA_X1 _3739_ (.A(_1721_),
    .B(_1722_),
    .CO(_1723_),
    .S(_1724_));
 HA_X1 _3740_ (.A(_1723_),
    .B(_1725_),
    .CO(_1726_),
    .S(_1727_));
 HA_X1 _3741_ (.A(_1728_),
    .B(_1729_),
    .CO(_1730_),
    .S(_1731_));
 HA_X1 _3742_ (.A(_1732_),
    .B(_1733_),
    .CO(_1734_),
    .S(_1735_));
 HA_X1 _3743_ (.A(_1736_),
    .B(_1737_),
    .CO(_1738_),
    .S(_1739_));
 HA_X1 _3744_ (.A(_1740_),
    .B(_1741_),
    .CO(_1742_),
    .S(_1743_));
 HA_X1 _3745_ (.A(_1744_),
    .B(_1745_),
    .CO(_1746_),
    .S(_1747_));
 HA_X1 _3746_ (.A(_1748_),
    .B(_1749_),
    .CO(_1750_),
    .S(_1751_));
 HA_X1 _3747_ (.A(_1752_),
    .B(_1753_),
    .CO(_1754_),
    .S(_1755_));
 HA_X1 _3748_ (.A(_1756_),
    .B(_1757_),
    .CO(_1758_),
    .S(_1759_));
 HA_X1 _3749_ (.A(_1760_),
    .B(_1761_),
    .CO(_1762_),
    .S(_1763_));
 HA_X1 _3750_ (.A(_1764_),
    .B(_1765_),
    .CO(_1766_),
    .S(_1767_));
 HA_X1 _3751_ (.A(_1768_),
    .B(net40),
    .CO(_1769_),
    .S(_1770_));
 HA_X1 _3752_ (.A(_1539_),
    .B(_1540_),
    .CO(_1771_),
    .S(_1772_));
 HA_X1 _3753_ (.A(net38),
    .B(_1535_),
    .CO(_1773_),
    .S(_1774_));
 HA_X1 _3754_ (.A(_1775_),
    .B(_1540_),
    .CO(_1776_),
    .S(_1777_));
 HA_X1 _3755_ (.A(net37),
    .B(_1535_),
    .CO(_1778_),
    .S(_1779_));
 HA_X1 _3756_ (.A(_1526_),
    .B(_1527_),
    .CO(_1780_),
    .S(_1781_));
 HA_X1 _3757_ (.A(net36),
    .B(_1531_),
    .CO(_1782_),
    .S(_1783_));
 HA_X1 _3758_ (.A(_1784_),
    .B(_1785_),
    .CO(_1786_),
    .S(_1787_));
 HA_X1 _3759_ (.A(net35),
    .B(_1788_),
    .CO(_1789_),
    .S(_1790_));
 HA_X1 _3760_ (.A(_1791_),
    .B(_1792_),
    .CO(_1793_),
    .S(_1794_));
 HA_X1 _3761_ (.A(_1522_),
    .B(_1523_),
    .CO(_1795_),
    .S(_1796_));
 HA_X1 _3762_ (.A(net34),
    .B(_1519_),
    .CO(_1797_),
    .S(_1798_));
 HA_X1 _3763_ (.A(_1799_),
    .B(_1800_),
    .CO(_1801_),
    .S(_1802_));
 HA_X1 _3764_ (.A(_1803_),
    .B(_1804_),
    .CO(_1791_),
    .S(_1805_));
 HA_X1 _3765_ (.A(_1806_),
    .B(_1807_),
    .CO(_1808_),
    .S(_1809_));
 HA_X1 _3766_ (.A(_1810_),
    .B(_1801_),
    .CO(_1811_),
    .S(_1812_));
 HA_X1 _3767_ (.A(net31),
    .B(_1813_),
    .CO(_1814_),
    .S(_1815_));
 HA_X1 _3768_ (.A(net30),
    .B(_1816_),
    .CO(_1817_),
    .S(_1818_));
 HA_X1 _3769_ (.A(net29),
    .B(_1819_),
    .CO(_1820_),
    .S(_1821_));
 HA_X1 _3770_ (.A(net27),
    .B(_1822_),
    .CO(_1823_),
    .S(_1824_));
 HA_X1 _3771_ (.A(net26),
    .B(_1825_),
    .CO(_1826_),
    .S(_1827_));
 HA_X1 _3772_ (.A(net25),
    .B(_1828_),
    .CO(_1829_),
    .S(_1830_));
 HA_X1 _3773_ (.A(net24),
    .B(_1831_),
    .CO(_1832_),
    .S(_1833_));
 HA_X1 _3774_ (.A(net23),
    .B(_1834_),
    .CO(_1835_),
    .S(_1836_));
 HA_X1 _3775_ (.A(net22),
    .B(_1837_),
    .CO(_1838_),
    .S(_1839_));
 HA_X1 _3776_ (.A(_1840_),
    .B(_1841_),
    .CO(_1516_),
    .S(_1842_));
 HA_X1 _3777_ (.A(net32),
    .B(_1843_),
    .CO(_1510_),
    .S(_1844_));
 HA_X1 _3778_ (.A(_1845_),
    .B(_1846_),
    .CO(_1847_),
    .S(_1848_));
 HA_X1 _3779_ (.A(_1550_),
    .B(_1551_),
    .CO(_1849_),
    .S(_1850_));
 HA_X1 _3780_ (.A(_1851_),
    .B(_1852_),
    .CO(_1853_),
    .S(_1854_));
 HA_X1 _3781_ (.A(_1555_),
    .B(_1556_),
    .CO(_1855_),
    .S(_1856_));
 HA_X1 _3782_ (.A(_1857_),
    .B(_1858_),
    .CO(_1859_),
    .S(_1860_));
 HA_X1 _3783_ (.A(_1560_),
    .B(_1561_),
    .CO(_1861_),
    .S(_1862_));
 HA_X1 _3784_ (.A(_1863_),
    .B(_1864_),
    .CO(_1865_),
    .S(_1866_));
 HA_X1 _3785_ (.A(_1565_),
    .B(_1566_),
    .CO(_1867_),
    .S(_1868_));
 HA_X1 _3786_ (.A(_1869_),
    .B(_1870_),
    .CO(_1871_),
    .S(_1872_));
 HA_X1 _3787_ (.A(_1873_),
    .B(_1874_),
    .CO(_1875_),
    .S(_1876_));
 HA_X1 _3788_ (.A(_1877_),
    .B(_1878_),
    .CO(_1879_),
    .S(_1880_));
 HA_X1 _3789_ (.A(_1575_),
    .B(_1576_),
    .CO(_1881_),
    .S(_1882_));
 HA_X1 _3790_ (.A(_1883_),
    .B(_1884_),
    .CO(_1885_),
    .S(_1886_));
 HA_X1 _3791_ (.A(_1887_),
    .B(_1888_),
    .CO(_1889_),
    .S(_1890_));
 HA_X1 _3792_ (.A(_1891_),
    .B(_1892_),
    .CO(_1893_),
    .S(_1894_));
 HA_X1 _3793_ (.A(_1895_),
    .B(_1896_),
    .CO(_1897_),
    .S(_1898_));
 HA_X1 _3794_ (.A(_1899_),
    .B(_1900_),
    .CO(_1901_),
    .S(_1902_));
 HA_X1 _3795_ (.A(_1903_),
    .B(_1904_),
    .CO(_1905_),
    .S(_1906_));
 HA_X1 _3796_ (.A(_1907_),
    .B(_1908_),
    .CO(_1909_),
    .S(_1910_));
 HA_X1 _3797_ (.A(_1911_),
    .B(_1912_),
    .CO(_1913_),
    .S(_1914_));
 HA_X1 _3798_ (.A(_1915_),
    .B(_1916_),
    .CO(_1917_),
    .S(_1918_));
 HA_X1 _3799_ (.A(_1919_),
    .B(_1920_),
    .CO(_1921_),
    .S(_1922_));
 HA_X1 _3800_ (.A(_1923_),
    .B(_1924_),
    .CO(_1925_),
    .S(_1926_));
 HA_X1 _3801_ (.A(_1605_),
    .B(_1222_),
    .CO(_1927_),
    .S(_1928_));
 HA_X1 _3802_ (.A(_1929_),
    .B(_1930_),
    .CO(_1931_),
    .S(_1932_));
 HA_X1 _3803_ (.A(_1196_),
    .B(_1134_),
    .CO(_1935_),
    .S(_1936_));
 HA_X1 _3804_ (.A(net97),
    .B(_1134_),
    .CO(_1937_),
    .S(_1938_));
 HA_X1 _3805_ (.A(_1842_),
    .B(_1135_),
    .CO(_1940_),
    .S(_1941_));
 HA_X1 _3806_ (.A(_1139_),
    .B(_1943_),
    .CO(_1944_),
    .S(_1945_));
 HA_X1 _3807_ (.A(_1946_),
    .B(_1947_),
    .CO(_1948_),
    .S(_1949_));
 TAPCELL_X1 PHY_0 ();
 BUF_X2 input42 (.A(operand_fp32_i[3]),
    .Z(net42));
 CLKBUF_X2 input43 (.A(operand_fp32_i[4]),
    .Z(net43));
 BUF_X2 input44 (.A(operand_fp32_i[5]),
    .Z(net44));
 BUF_X2 input45 (.A(operand_fp32_i[6]),
    .Z(net45));
 BUF_X2 input46 (.A(operand_fp32_i[7]),
    .Z(net46));
 BUF_X2 input47 (.A(operand_fp32_i[8]),
    .Z(net47));
 BUF_X2 input48 (.A(operand_fp32_i[9]),
    .Z(net48));
 BUF_X4 output49 (.A(net49),
    .Z(result_o[0]));
 BUF_X4 output50 (.A(net50),
    .Z(result_o[10]));
 BUF_X4 output51 (.A(net51),
    .Z(result_o[11]));
 BUF_X4 output52 (.A(net52),
    .Z(result_o[12]));
 BUF_X4 output53 (.A(net53),
    .Z(result_o[13]));
 BUF_X4 output54 (.A(net54),
    .Z(result_o[14]));
 BUF_X4 output55 (.A(net55),
    .Z(result_o[15]));
 BUF_X4 output56 (.A(net56),
    .Z(result_o[16]));
 BUF_X4 output57 (.A(net57),
    .Z(result_o[17]));
 BUF_X4 output58 (.A(net58),
    .Z(result_o[18]));
 BUF_X4 output59 (.A(net59),
    .Z(result_o[19]));
 BUF_X4 output60 (.A(net60),
    .Z(result_o[1]));
 BUF_X4 output61 (.A(net61),
    .Z(result_o[20]));
 BUF_X4 output62 (.A(net62),
    .Z(result_o[21]));
 BUF_X4 output63 (.A(net63),
    .Z(result_o[22]));
 BUF_X4 output64 (.A(net64),
    .Z(result_o[23]));
 BUF_X4 output65 (.A(net65),
    .Z(result_o[24]));
 BUF_X4 output66 (.A(net66),
    .Z(result_o[25]));
 BUF_X4 output67 (.A(net67),
    .Z(result_o[26]));
 BUF_X4 output68 (.A(net68),
    .Z(result_o[27]));
 BUF_X4 output69 (.A(net69),
    .Z(result_o[28]));
 BUF_X4 output70 (.A(net70),
    .Z(result_o[29]));
 BUF_X4 output71 (.A(net71),
    .Z(result_o[2]));
 BUF_X4 output72 (.A(net72),
    .Z(result_o[30]));
 BUF_X4 output73 (.A(net73),
    .Z(result_o[31]));
 BUF_X4 output74 (.A(net74),
    .Z(result_o[3]));
 BUF_X4 output75 (.A(net75),
    .Z(result_o[4]));
 BUF_X4 output76 (.A(net76),
    .Z(result_o[5]));
 BUF_X4 output77 (.A(net77),
    .Z(result_o[6]));
 BUF_X4 output78 (.A(net78),
    .Z(result_o[7]));
 BUF_X4 output79 (.A(net79),
    .Z(result_o[8]));
 BUF_X4 output80 (.A(net80),
    .Z(result_o[9]));
 BUF_X4 max_cap81 (.A(_0737_),
    .Z(net81));
 BUF_X8 wire82 (.A(_1700_),
    .Z(net82));
 BUF_X4 max_cap83 (.A(_1693_),
    .Z(net83));
 BUF_X4 max_cap84 (.A(net85),
    .Z(net84));
 BUF_X4 max_cap85 (.A(_1687_),
    .Z(net85));
 BUF_X16 max_cap86 (.A(_0117_),
    .Z(net86));
 BUF_X4 max_cap87 (.A(_1681_),
    .Z(net87));
 BUF_X2 max_cap88 (.A(_1945_),
    .Z(net88));
 BUF_X4 max_cap89 (.A(_1936_),
    .Z(net89));
 BUF_X4 max_cap90 (.A(net92),
    .Z(net90));
 BUF_X4 max_cap91 (.A(net92),
    .Z(net91));
 BUF_X4 max_cap92 (.A(_1123_),
    .Z(net92));
 CLKBUF_X3 wire93 (.A(net96),
    .Z(net93));
 BUF_X4 max_cap94 (.A(net95),
    .Z(net94));
 CLKBUF_X3 max_cap95 (.A(net97),
    .Z(net95));
 BUF_X4 max_cap96 (.A(net97),
    .Z(net96));
 CLKBUF_X3 max_cap97 (.A(_1842_),
    .Z(net97));
 BUF_X4 max_cap98 (.A(_1802_),
    .Z(net98));
 FILLCELL_X32 FILLER_0_0_1 ();
 FILLCELL_X32 FILLER_0_0_33 ();
 FILLCELL_X16 FILLER_0_0_65 ();
 FILLCELL_X4 FILLER_0_0_81 ();
 FILLCELL_X2 FILLER_0_0_85 ();
 FILLCELL_X4 FILLER_0_0_92 ();
 FILLCELL_X2 FILLER_0_0_96 ();
 FILLCELL_X8 FILLER_0_0_102 ();
 FILLCELL_X32 FILLER_0_0_113 ();
 FILLCELL_X2 FILLER_0_0_149 ();
 FILLCELL_X1 FILLER_0_0_151 ();
 FILLCELL_X16 FILLER_0_0_159 ();
 FILLCELL_X8 FILLER_0_0_175 ();
 FILLCELL_X4 FILLER_0_0_183 ();
 FILLCELL_X8 FILLER_0_0_194 ();
 FILLCELL_X4 FILLER_0_0_209 ();
 FILLCELL_X1 FILLER_0_0_213 ();
 FILLCELL_X8 FILLER_0_0_228 ();
 FILLCELL_X2 FILLER_0_0_236 ();
 FILLCELL_X8 FILLER_0_0_247 ();
 FILLCELL_X2 FILLER_0_0_255 ();
 FILLCELL_X32 FILLER_0_0_264 ();
 FILLCELL_X32 FILLER_0_0_296 ();
 FILLCELL_X32 FILLER_0_0_328 ();
 FILLCELL_X32 FILLER_0_0_360 ();
 FILLCELL_X16 FILLER_0_0_392 ();
 FILLCELL_X2 FILLER_0_0_408 ();
 FILLCELL_X1 FILLER_0_0_410 ();
 FILLCELL_X32 FILLER_0_1_1 ();
 FILLCELL_X32 FILLER_0_1_33 ();
 FILLCELL_X32 FILLER_0_1_65 ();
 FILLCELL_X32 FILLER_0_1_97 ();
 FILLCELL_X8 FILLER_0_1_129 ();
 FILLCELL_X2 FILLER_0_1_137 ();
 FILLCELL_X32 FILLER_0_1_142 ();
 FILLCELL_X16 FILLER_0_1_174 ();
 FILLCELL_X4 FILLER_0_1_190 ();
 FILLCELL_X1 FILLER_0_1_194 ();
 FILLCELL_X32 FILLER_0_1_204 ();
 FILLCELL_X16 FILLER_0_1_236 ();
 FILLCELL_X4 FILLER_0_1_252 ();
 FILLCELL_X2 FILLER_0_1_256 ();
 FILLCELL_X1 FILLER_0_1_260 ();
 FILLCELL_X32 FILLER_0_1_268 ();
 FILLCELL_X32 FILLER_0_1_300 ();
 FILLCELL_X32 FILLER_0_1_332 ();
 FILLCELL_X32 FILLER_0_1_364 ();
 FILLCELL_X8 FILLER_0_1_396 ();
 FILLCELL_X4 FILLER_0_1_404 ();
 FILLCELL_X2 FILLER_0_1_408 ();
 FILLCELL_X1 FILLER_0_1_410 ();
 FILLCELL_X32 FILLER_0_2_1 ();
 FILLCELL_X32 FILLER_0_2_33 ();
 FILLCELL_X32 FILLER_0_2_65 ();
 FILLCELL_X32 FILLER_0_2_97 ();
 FILLCELL_X32 FILLER_0_2_129 ();
 FILLCELL_X32 FILLER_0_2_161 ();
 FILLCELL_X32 FILLER_0_2_193 ();
 FILLCELL_X32 FILLER_0_2_225 ();
 FILLCELL_X32 FILLER_0_2_257 ();
 FILLCELL_X32 FILLER_0_2_289 ();
 FILLCELL_X32 FILLER_0_2_321 ();
 FILLCELL_X32 FILLER_0_2_353 ();
 FILLCELL_X16 FILLER_0_2_385 ();
 FILLCELL_X8 FILLER_0_2_401 ();
 FILLCELL_X2 FILLER_0_2_409 ();
 FILLCELL_X32 FILLER_0_3_1 ();
 FILLCELL_X32 FILLER_0_3_33 ();
 FILLCELL_X32 FILLER_0_3_65 ();
 FILLCELL_X32 FILLER_0_3_97 ();
 FILLCELL_X32 FILLER_0_3_129 ();
 FILLCELL_X32 FILLER_0_3_161 ();
 FILLCELL_X8 FILLER_0_3_193 ();
 FILLCELL_X1 FILLER_0_3_201 ();
 FILLCELL_X16 FILLER_0_3_209 ();
 FILLCELL_X8 FILLER_0_3_225 ();
 FILLCELL_X32 FILLER_0_3_243 ();
 FILLCELL_X32 FILLER_0_3_275 ();
 FILLCELL_X32 FILLER_0_3_307 ();
 FILLCELL_X32 FILLER_0_3_339 ();
 FILLCELL_X32 FILLER_0_3_371 ();
 FILLCELL_X8 FILLER_0_3_403 ();
 FILLCELL_X32 FILLER_0_4_1 ();
 FILLCELL_X32 FILLER_0_4_33 ();
 FILLCELL_X32 FILLER_0_4_65 ();
 FILLCELL_X32 FILLER_0_4_97 ();
 FILLCELL_X8 FILLER_0_4_129 ();
 FILLCELL_X32 FILLER_0_4_139 ();
 FILLCELL_X16 FILLER_0_4_171 ();
 FILLCELL_X8 FILLER_0_4_187 ();
 FILLCELL_X2 FILLER_0_4_247 ();
 FILLCELL_X32 FILLER_0_4_251 ();
 FILLCELL_X32 FILLER_0_4_283 ();
 FILLCELL_X32 FILLER_0_4_315 ();
 FILLCELL_X32 FILLER_0_4_347 ();
 FILLCELL_X32 FILLER_0_4_379 ();
 FILLCELL_X16 FILLER_0_5_1 ();
 FILLCELL_X8 FILLER_0_5_17 ();
 FILLCELL_X4 FILLER_0_5_25 ();
 FILLCELL_X2 FILLER_0_5_29 ();
 FILLCELL_X32 FILLER_0_5_37 ();
 FILLCELL_X16 FILLER_0_5_69 ();
 FILLCELL_X8 FILLER_0_5_85 ();
 FILLCELL_X2 FILLER_0_5_117 ();
 FILLCELL_X8 FILLER_0_5_123 ();
 FILLCELL_X4 FILLER_0_5_131 ();
 FILLCELL_X32 FILLER_0_5_145 ();
 FILLCELL_X4 FILLER_0_5_177 ();
 FILLCELL_X1 FILLER_0_5_181 ();
 FILLCELL_X1 FILLER_0_5_204 ();
 FILLCELL_X1 FILLER_0_5_215 ();
 FILLCELL_X8 FILLER_0_5_230 ();
 FILLCELL_X1 FILLER_0_5_238 ();
 FILLCELL_X32 FILLER_0_5_261 ();
 FILLCELL_X32 FILLER_0_5_293 ();
 FILLCELL_X32 FILLER_0_5_325 ();
 FILLCELL_X32 FILLER_0_5_357 ();
 FILLCELL_X16 FILLER_0_5_389 ();
 FILLCELL_X4 FILLER_0_5_405 ();
 FILLCELL_X2 FILLER_0_5_409 ();
 FILLCELL_X4 FILLER_0_6_1 ();
 FILLCELL_X8 FILLER_0_6_7 ();
 FILLCELL_X4 FILLER_0_6_15 ();
 FILLCELL_X1 FILLER_0_6_21 ();
 FILLCELL_X1 FILLER_0_6_26 ();
 FILLCELL_X1 FILLER_0_6_31 ();
 FILLCELL_X1 FILLER_0_6_40 ();
 FILLCELL_X32 FILLER_0_6_48 ();
 FILLCELL_X8 FILLER_0_6_80 ();
 FILLCELL_X2 FILLER_0_6_88 ();
 FILLCELL_X2 FILLER_0_6_112 ();
 FILLCELL_X1 FILLER_0_6_143 ();
 FILLCELL_X4 FILLER_0_6_148 ();
 FILLCELL_X2 FILLER_0_6_152 ();
 FILLCELL_X1 FILLER_0_6_154 ();
 FILLCELL_X32 FILLER_0_6_165 ();
 FILLCELL_X2 FILLER_0_6_197 ();
 FILLCELL_X2 FILLER_0_6_206 ();
 FILLCELL_X8 FILLER_0_6_210 ();
 FILLCELL_X1 FILLER_0_6_218 ();
 FILLCELL_X2 FILLER_0_6_223 ();
 FILLCELL_X4 FILLER_0_6_229 ();
 FILLCELL_X1 FILLER_0_6_233 ();
 FILLCELL_X4 FILLER_0_6_256 ();
 FILLCELL_X32 FILLER_0_6_270 ();
 FILLCELL_X32 FILLER_0_6_302 ();
 FILLCELL_X32 FILLER_0_6_334 ();
 FILLCELL_X32 FILLER_0_6_366 ();
 FILLCELL_X8 FILLER_0_6_398 ();
 FILLCELL_X4 FILLER_0_6_406 ();
 FILLCELL_X1 FILLER_0_6_410 ();
 FILLCELL_X2 FILLER_0_7_14 ();
 FILLCELL_X1 FILLER_0_7_46 ();
 FILLCELL_X2 FILLER_0_7_54 ();
 FILLCELL_X1 FILLER_0_7_56 ();
 FILLCELL_X8 FILLER_0_7_67 ();
 FILLCELL_X4 FILLER_0_7_75 ();
 FILLCELL_X2 FILLER_0_7_79 ();
 FILLCELL_X1 FILLER_0_7_113 ();
 FILLCELL_X2 FILLER_0_7_164 ();
 FILLCELL_X8 FILLER_0_7_175 ();
 FILLCELL_X4 FILLER_0_7_183 ();
 FILLCELL_X4 FILLER_0_7_199 ();
 FILLCELL_X2 FILLER_0_7_213 ();
 FILLCELL_X32 FILLER_0_7_269 ();
 FILLCELL_X32 FILLER_0_7_301 ();
 FILLCELL_X32 FILLER_0_7_333 ();
 FILLCELL_X32 FILLER_0_7_365 ();
 FILLCELL_X8 FILLER_0_7_397 ();
 FILLCELL_X4 FILLER_0_7_405 ();
 FILLCELL_X2 FILLER_0_7_409 ();
 FILLCELL_X1 FILLER_0_8_1 ();
 FILLCELL_X1 FILLER_0_8_15 ();
 FILLCELL_X1 FILLER_0_8_19 ();
 FILLCELL_X1 FILLER_0_8_23 ();
 FILLCELL_X1 FILLER_0_8_37 ();
 FILLCELL_X2 FILLER_0_8_56 ();
 FILLCELL_X1 FILLER_0_8_58 ();
 FILLCELL_X2 FILLER_0_8_61 ();
 FILLCELL_X1 FILLER_0_8_63 ();
 FILLCELL_X1 FILLER_0_8_77 ();
 FILLCELL_X1 FILLER_0_8_81 ();
 FILLCELL_X4 FILLER_0_8_91 ();
 FILLCELL_X2 FILLER_0_8_95 ();
 FILLCELL_X1 FILLER_0_8_112 ();
 FILLCELL_X1 FILLER_0_8_121 ();
 FILLCELL_X1 FILLER_0_8_124 ();
 FILLCELL_X1 FILLER_0_8_129 ();
 FILLCELL_X4 FILLER_0_8_143 ();
 FILLCELL_X2 FILLER_0_8_153 ();
 FILLCELL_X16 FILLER_0_8_178 ();
 FILLCELL_X4 FILLER_0_8_196 ();
 FILLCELL_X2 FILLER_0_8_200 ();
 FILLCELL_X1 FILLER_0_8_212 ();
 FILLCELL_X4 FILLER_0_8_223 ();
 FILLCELL_X1 FILLER_0_8_227 ();
 FILLCELL_X4 FILLER_0_8_254 ();
 FILLCELL_X2 FILLER_0_8_258 ();
 FILLCELL_X4 FILLER_0_8_265 ();
 FILLCELL_X1 FILLER_0_8_269 ();
 FILLCELL_X16 FILLER_0_8_275 ();
 FILLCELL_X8 FILLER_0_8_301 ();
 FILLCELL_X32 FILLER_0_8_315 ();
 FILLCELL_X32 FILLER_0_8_347 ();
 FILLCELL_X32 FILLER_0_8_379 ();
 FILLCELL_X1 FILLER_0_9_26 ();
 FILLCELL_X1 FILLER_0_9_29 ();
 FILLCELL_X1 FILLER_0_9_35 ();
 FILLCELL_X1 FILLER_0_9_39 ();
 FILLCELL_X1 FILLER_0_9_61 ();
 FILLCELL_X1 FILLER_0_9_72 ();
 FILLCELL_X1 FILLER_0_9_80 ();
 FILLCELL_X2 FILLER_0_9_94 ();
 FILLCELL_X4 FILLER_0_9_122 ();
 FILLCELL_X2 FILLER_0_9_126 ();
 FILLCELL_X1 FILLER_0_9_128 ();
 FILLCELL_X2 FILLER_0_9_155 ();
 FILLCELL_X16 FILLER_0_9_174 ();
 FILLCELL_X8 FILLER_0_9_190 ();
 FILLCELL_X2 FILLER_0_9_198 ();
 FILLCELL_X1 FILLER_0_9_200 ();
 FILLCELL_X2 FILLER_0_9_213 ();
 FILLCELL_X4 FILLER_0_9_244 ();
 FILLCELL_X2 FILLER_0_9_248 ();
 FILLCELL_X1 FILLER_0_9_255 ();
 FILLCELL_X2 FILLER_0_9_269 ();
 FILLCELL_X8 FILLER_0_9_284 ();
 FILLCELL_X1 FILLER_0_9_292 ();
 FILLCELL_X2 FILLER_0_9_311 ();
 FILLCELL_X1 FILLER_0_9_313 ();
 FILLCELL_X32 FILLER_0_9_320 ();
 FILLCELL_X32 FILLER_0_9_352 ();
 FILLCELL_X16 FILLER_0_9_384 ();
 FILLCELL_X8 FILLER_0_9_400 ();
 FILLCELL_X2 FILLER_0_9_408 ();
 FILLCELL_X1 FILLER_0_9_410 ();
 FILLCELL_X1 FILLER_0_10_1 ();
 FILLCELL_X1 FILLER_0_10_59 ();
 FILLCELL_X1 FILLER_0_10_67 ();
 FILLCELL_X2 FILLER_0_10_73 ();
 FILLCELL_X1 FILLER_0_10_80 ();
 FILLCELL_X1 FILLER_0_10_94 ();
 FILLCELL_X1 FILLER_0_10_105 ();
 FILLCELL_X1 FILLER_0_10_108 ();
 FILLCELL_X4 FILLER_0_10_119 ();
 FILLCELL_X1 FILLER_0_10_143 ();
 FILLCELL_X16 FILLER_0_10_169 ();
 FILLCELL_X8 FILLER_0_10_185 ();
 FILLCELL_X4 FILLER_0_10_193 ();
 FILLCELL_X2 FILLER_0_10_197 ();
 FILLCELL_X1 FILLER_0_10_223 ();
 FILLCELL_X1 FILLER_0_10_230 ();
 FILLCELL_X1 FILLER_0_10_233 ();
 FILLCELL_X1 FILLER_0_10_236 ();
 FILLCELL_X1 FILLER_0_10_247 ();
 FILLCELL_X1 FILLER_0_10_268 ();
 FILLCELL_X8 FILLER_0_10_300 ();
 FILLCELL_X2 FILLER_0_10_314 ();
 FILLCELL_X32 FILLER_0_10_326 ();
 FILLCELL_X32 FILLER_0_10_358 ();
 FILLCELL_X16 FILLER_0_10_390 ();
 FILLCELL_X4 FILLER_0_10_406 ();
 FILLCELL_X1 FILLER_0_10_410 ();
 FILLCELL_X2 FILLER_0_11_47 ();
 FILLCELL_X8 FILLER_0_11_53 ();
 FILLCELL_X4 FILLER_0_11_61 ();
 FILLCELL_X1 FILLER_0_11_65 ();
 FILLCELL_X8 FILLER_0_11_89 ();
 FILLCELL_X2 FILLER_0_11_97 ();
 FILLCELL_X1 FILLER_0_11_99 ();
 FILLCELL_X4 FILLER_0_11_108 ();
 FILLCELL_X2 FILLER_0_11_112 ();
 FILLCELL_X4 FILLER_0_11_123 ();
 FILLCELL_X2 FILLER_0_11_127 ();
 FILLCELL_X1 FILLER_0_11_129 ();
 FILLCELL_X4 FILLER_0_11_146 ();
 FILLCELL_X32 FILLER_0_11_166 ();
 FILLCELL_X4 FILLER_0_11_198 ();
 FILLCELL_X2 FILLER_0_11_202 ();
 FILLCELL_X1 FILLER_0_11_204 ();
 FILLCELL_X16 FILLER_0_11_207 ();
 FILLCELL_X2 FILLER_0_11_223 ();
 FILLCELL_X1 FILLER_0_11_225 ();
 FILLCELL_X16 FILLER_0_11_239 ();
 FILLCELL_X4 FILLER_0_11_255 ();
 FILLCELL_X2 FILLER_0_11_259 ();
 FILLCELL_X1 FILLER_0_11_261 ();
 FILLCELL_X2 FILLER_0_11_273 ();
 FILLCELL_X1 FILLER_0_11_275 ();
 FILLCELL_X2 FILLER_0_11_287 ();
 FILLCELL_X1 FILLER_0_11_315 ();
 FILLCELL_X32 FILLER_0_11_338 ();
 FILLCELL_X32 FILLER_0_11_370 ();
 FILLCELL_X8 FILLER_0_11_402 ();
 FILLCELL_X1 FILLER_0_11_410 ();
 FILLCELL_X2 FILLER_0_12_97 ();
 FILLCELL_X4 FILLER_0_12_119 ();
 FILLCELL_X2 FILLER_0_12_123 ();
 FILLCELL_X1 FILLER_0_12_125 ();
 FILLCELL_X2 FILLER_0_12_135 ();
 FILLCELL_X1 FILLER_0_12_137 ();
 FILLCELL_X8 FILLER_0_12_156 ();
 FILLCELL_X1 FILLER_0_12_164 ();
 FILLCELL_X16 FILLER_0_12_174 ();
 FILLCELL_X4 FILLER_0_12_190 ();
 FILLCELL_X2 FILLER_0_12_194 ();
 FILLCELL_X1 FILLER_0_12_196 ();
 FILLCELL_X4 FILLER_0_12_209 ();
 FILLCELL_X2 FILLER_0_12_213 ();
 FILLCELL_X1 FILLER_0_12_215 ();
 FILLCELL_X2 FILLER_0_12_224 ();
 FILLCELL_X2 FILLER_0_12_242 ();
 FILLCELL_X1 FILLER_0_12_244 ();
 FILLCELL_X1 FILLER_0_12_274 ();
 FILLCELL_X4 FILLER_0_12_298 ();
 FILLCELL_X2 FILLER_0_12_302 ();
 FILLCELL_X1 FILLER_0_12_304 ();
 FILLCELL_X1 FILLER_0_12_309 ();
 FILLCELL_X1 FILLER_0_12_321 ();
 FILLCELL_X2 FILLER_0_12_326 ();
 FILLCELL_X32 FILLER_0_12_345 ();
 FILLCELL_X32 FILLER_0_12_377 ();
 FILLCELL_X2 FILLER_0_12_409 ();
 FILLCELL_X2 FILLER_0_13_67 ();
 FILLCELL_X1 FILLER_0_13_73 ();
 FILLCELL_X2 FILLER_0_13_81 ();
 FILLCELL_X1 FILLER_0_13_83 ();
 FILLCELL_X2 FILLER_0_13_121 ();
 FILLCELL_X8 FILLER_0_13_142 ();
 FILLCELL_X1 FILLER_0_13_150 ();
 FILLCELL_X32 FILLER_0_13_161 ();
 FILLCELL_X2 FILLER_0_13_193 ();
 FILLCELL_X2 FILLER_0_13_213 ();
 FILLCELL_X1 FILLER_0_13_215 ();
 FILLCELL_X1 FILLER_0_13_219 ();
 FILLCELL_X2 FILLER_0_13_225 ();
 FILLCELL_X2 FILLER_0_13_232 ();
 FILLCELL_X1 FILLER_0_13_234 ();
 FILLCELL_X4 FILLER_0_13_260 ();
 FILLCELL_X1 FILLER_0_13_264 ();
 FILLCELL_X1 FILLER_0_13_271 ();
 FILLCELL_X2 FILLER_0_13_279 ();
 FILLCELL_X1 FILLER_0_13_283 ();
 FILLCELL_X1 FILLER_0_13_296 ();
 FILLCELL_X2 FILLER_0_13_300 ();
 FILLCELL_X32 FILLER_0_13_341 ();
 FILLCELL_X32 FILLER_0_13_373 ();
 FILLCELL_X4 FILLER_0_13_405 ();
 FILLCELL_X2 FILLER_0_13_409 ();
 FILLCELL_X1 FILLER_0_14_32 ();
 FILLCELL_X8 FILLER_0_14_56 ();
 FILLCELL_X1 FILLER_0_14_64 ();
 FILLCELL_X2 FILLER_0_14_75 ();
 FILLCELL_X1 FILLER_0_14_77 ();
 FILLCELL_X8 FILLER_0_14_85 ();
 FILLCELL_X4 FILLER_0_14_93 ();
 FILLCELL_X2 FILLER_0_14_113 ();
 FILLCELL_X1 FILLER_0_14_115 ();
 FILLCELL_X2 FILLER_0_14_122 ();
 FILLCELL_X4 FILLER_0_14_143 ();
 FILLCELL_X2 FILLER_0_14_147 ();
 FILLCELL_X2 FILLER_0_14_153 ();
 FILLCELL_X2 FILLER_0_14_192 ();
 FILLCELL_X1 FILLER_0_14_198 ();
 FILLCELL_X2 FILLER_0_14_203 ();
 FILLCELL_X1 FILLER_0_14_216 ();
 FILLCELL_X4 FILLER_0_14_229 ();
 FILLCELL_X2 FILLER_0_14_233 ();
 FILLCELL_X4 FILLER_0_14_238 ();
 FILLCELL_X1 FILLER_0_14_242 ();
 FILLCELL_X2 FILLER_0_14_256 ();
 FILLCELL_X2 FILLER_0_14_267 ();
 FILLCELL_X1 FILLER_0_14_269 ();
 FILLCELL_X4 FILLER_0_14_305 ();
 FILLCELL_X2 FILLER_0_14_309 ();
 FILLCELL_X1 FILLER_0_14_311 ();
 FILLCELL_X32 FILLER_0_14_342 ();
 FILLCELL_X32 FILLER_0_14_374 ();
 FILLCELL_X4 FILLER_0_14_406 ();
 FILLCELL_X1 FILLER_0_14_410 ();
 FILLCELL_X4 FILLER_0_15_56 ();
 FILLCELL_X2 FILLER_0_15_60 ();
 FILLCELL_X2 FILLER_0_15_70 ();
 FILLCELL_X1 FILLER_0_15_72 ();
 FILLCELL_X2 FILLER_0_15_80 ();
 FILLCELL_X1 FILLER_0_15_82 ();
 FILLCELL_X1 FILLER_0_15_87 ();
 FILLCELL_X1 FILLER_0_15_98 ();
 FILLCELL_X2 FILLER_0_15_102 ();
 FILLCELL_X1 FILLER_0_15_104 ();
 FILLCELL_X1 FILLER_0_15_112 ();
 FILLCELL_X8 FILLER_0_15_122 ();
 FILLCELL_X2 FILLER_0_15_130 ();
 FILLCELL_X4 FILLER_0_15_144 ();
 FILLCELL_X1 FILLER_0_15_148 ();
 FILLCELL_X4 FILLER_0_15_165 ();
 FILLCELL_X1 FILLER_0_15_169 ();
 FILLCELL_X1 FILLER_0_15_180 ();
 FILLCELL_X1 FILLER_0_15_198 ();
 FILLCELL_X1 FILLER_0_15_206 ();
 FILLCELL_X1 FILLER_0_15_211 ();
 FILLCELL_X2 FILLER_0_15_221 ();
 FILLCELL_X1 FILLER_0_15_240 ();
 FILLCELL_X2 FILLER_0_15_250 ();
 FILLCELL_X1 FILLER_0_15_268 ();
 FILLCELL_X1 FILLER_0_15_302 ();
 FILLCELL_X4 FILLER_0_15_332 ();
 FILLCELL_X2 FILLER_0_15_336 ();
 FILLCELL_X1 FILLER_0_15_338 ();
 FILLCELL_X32 FILLER_0_15_352 ();
 FILLCELL_X16 FILLER_0_15_384 ();
 FILLCELL_X8 FILLER_0_15_400 ();
 FILLCELL_X2 FILLER_0_15_408 ();
 FILLCELL_X1 FILLER_0_15_410 ();
 FILLCELL_X1 FILLER_0_16_31 ();
 FILLCELL_X2 FILLER_0_16_50 ();
 FILLCELL_X1 FILLER_0_16_70 ();
 FILLCELL_X4 FILLER_0_16_95 ();
 FILLCELL_X8 FILLER_0_16_106 ();
 FILLCELL_X1 FILLER_0_16_114 ();
 FILLCELL_X1 FILLER_0_16_121 ();
 FILLCELL_X4 FILLER_0_16_132 ();
 FILLCELL_X2 FILLER_0_16_136 ();
 FILLCELL_X1 FILLER_0_16_138 ();
 FILLCELL_X16 FILLER_0_16_159 ();
 FILLCELL_X4 FILLER_0_16_175 ();
 FILLCELL_X1 FILLER_0_16_179 ();
 FILLCELL_X4 FILLER_0_16_184 ();
 FILLCELL_X2 FILLER_0_16_188 ();
 FILLCELL_X2 FILLER_0_16_206 ();
 FILLCELL_X1 FILLER_0_16_228 ();
 FILLCELL_X4 FILLER_0_16_247 ();
 FILLCELL_X4 FILLER_0_16_258 ();
 FILLCELL_X4 FILLER_0_16_270 ();
 FILLCELL_X1 FILLER_0_16_274 ();
 FILLCELL_X2 FILLER_0_16_284 ();
 FILLCELL_X1 FILLER_0_16_293 ();
 FILLCELL_X1 FILLER_0_16_300 ();
 FILLCELL_X1 FILLER_0_16_310 ();
 FILLCELL_X2 FILLER_0_16_315 ();
 FILLCELL_X1 FILLER_0_16_317 ();
 FILLCELL_X1 FILLER_0_16_329 ();
 FILLCELL_X1 FILLER_0_16_333 ();
 FILLCELL_X1 FILLER_0_16_343 ();
 FILLCELL_X1 FILLER_0_16_348 ();
 FILLCELL_X1 FILLER_0_16_352 ();
 FILLCELL_X1 FILLER_0_16_359 ();
 FILLCELL_X1 FILLER_0_16_365 ();
 FILLCELL_X1 FILLER_0_16_369 ();
 FILLCELL_X1 FILLER_0_16_373 ();
 FILLCELL_X32 FILLER_0_16_379 ();
 FILLCELL_X8 FILLER_0_17_81 ();
 FILLCELL_X4 FILLER_0_17_89 ();
 FILLCELL_X1 FILLER_0_17_93 ();
 FILLCELL_X8 FILLER_0_17_96 ();
 FILLCELL_X2 FILLER_0_17_113 ();
 FILLCELL_X1 FILLER_0_17_115 ();
 FILLCELL_X1 FILLER_0_17_122 ();
 FILLCELL_X8 FILLER_0_17_159 ();
 FILLCELL_X4 FILLER_0_17_167 ();
 FILLCELL_X2 FILLER_0_17_171 ();
 FILLCELL_X8 FILLER_0_17_189 ();
 FILLCELL_X1 FILLER_0_17_202 ();
 FILLCELL_X8 FILLER_0_17_207 ();
 FILLCELL_X4 FILLER_0_17_215 ();
 FILLCELL_X2 FILLER_0_17_241 ();
 FILLCELL_X2 FILLER_0_17_251 ();
 FILLCELL_X1 FILLER_0_17_253 ();
 FILLCELL_X2 FILLER_0_17_298 ();
 FILLCELL_X1 FILLER_0_17_320 ();
 FILLCELL_X1 FILLER_0_17_352 ();
 FILLCELL_X4 FILLER_0_17_378 ();
 FILLCELL_X1 FILLER_0_17_382 ();
 FILLCELL_X8 FILLER_0_17_399 ();
 FILLCELL_X4 FILLER_0_17_407 ();
 FILLCELL_X2 FILLER_0_18_13 ();
 FILLCELL_X2 FILLER_0_18_63 ();
 FILLCELL_X1 FILLER_0_18_78 ();
 FILLCELL_X2 FILLER_0_18_88 ();
 FILLCELL_X2 FILLER_0_18_96 ();
 FILLCELL_X2 FILLER_0_18_112 ();
 FILLCELL_X2 FILLER_0_18_118 ();
 FILLCELL_X1 FILLER_0_18_120 ();
 FILLCELL_X2 FILLER_0_18_127 ();
 FILLCELL_X1 FILLER_0_18_129 ();
 FILLCELL_X2 FILLER_0_18_140 ();
 FILLCELL_X8 FILLER_0_18_164 ();
 FILLCELL_X1 FILLER_0_18_172 ();
 FILLCELL_X4 FILLER_0_18_220 ();
 FILLCELL_X2 FILLER_0_18_224 ();
 FILLCELL_X1 FILLER_0_18_226 ();
 FILLCELL_X4 FILLER_0_18_230 ();
 FILLCELL_X1 FILLER_0_18_234 ();
 FILLCELL_X4 FILLER_0_18_250 ();
 FILLCELL_X8 FILLER_0_18_261 ();
 FILLCELL_X4 FILLER_0_18_269 ();
 FILLCELL_X2 FILLER_0_18_273 ();
 FILLCELL_X4 FILLER_0_18_287 ();
 FILLCELL_X2 FILLER_0_18_291 ();
 FILLCELL_X1 FILLER_0_18_321 ();
 FILLCELL_X2 FILLER_0_18_347 ();
 FILLCELL_X8 FILLER_0_18_365 ();
 FILLCELL_X4 FILLER_0_18_373 ();
 FILLCELL_X2 FILLER_0_18_377 ();
 FILLCELL_X8 FILLER_0_18_384 ();
 FILLCELL_X1 FILLER_0_18_392 ();
 FILLCELL_X4 FILLER_0_18_406 ();
 FILLCELL_X1 FILLER_0_18_410 ();
 FILLCELL_X1 FILLER_0_19_28 ();
 FILLCELL_X1 FILLER_0_19_33 ();
 FILLCELL_X1 FILLER_0_19_38 ();
 FILLCELL_X1 FILLER_0_19_47 ();
 FILLCELL_X2 FILLER_0_19_51 ();
 FILLCELL_X1 FILLER_0_19_123 ();
 FILLCELL_X2 FILLER_0_19_130 ();
 FILLCELL_X1 FILLER_0_19_135 ();
 FILLCELL_X2 FILLER_0_19_145 ();
 FILLCELL_X8 FILLER_0_19_182 ();
 FILLCELL_X4 FILLER_0_19_190 ();
 FILLCELL_X4 FILLER_0_19_200 ();
 FILLCELL_X1 FILLER_0_19_204 ();
 FILLCELL_X4 FILLER_0_19_219 ();
 FILLCELL_X1 FILLER_0_19_223 ();
 FILLCELL_X4 FILLER_0_19_228 ();
 FILLCELL_X2 FILLER_0_19_232 ();
 FILLCELL_X4 FILLER_0_19_252 ();
 FILLCELL_X2 FILLER_0_19_256 ();
 FILLCELL_X4 FILLER_0_19_272 ();
 FILLCELL_X1 FILLER_0_19_276 ();
 FILLCELL_X8 FILLER_0_19_289 ();
 FILLCELL_X1 FILLER_0_19_297 ();
 FILLCELL_X1 FILLER_0_19_302 ();
 FILLCELL_X1 FILLER_0_19_329 ();
 FILLCELL_X2 FILLER_0_19_336 ();
 FILLCELL_X2 FILLER_0_19_354 ();
 FILLCELL_X4 FILLER_0_19_370 ();
 FILLCELL_X1 FILLER_0_19_374 ();
 FILLCELL_X2 FILLER_0_19_383 ();
 FILLCELL_X2 FILLER_0_19_402 ();
 FILLCELL_X1 FILLER_0_20_1 ();
 FILLCELL_X1 FILLER_0_20_42 ();
 FILLCELL_X1 FILLER_0_20_46 ();
 FILLCELL_X1 FILLER_0_20_57 ();
 FILLCELL_X1 FILLER_0_20_68 ();
 FILLCELL_X1 FILLER_0_20_73 ();
 FILLCELL_X1 FILLER_0_20_97 ();
 FILLCELL_X1 FILLER_0_20_104 ();
 FILLCELL_X4 FILLER_0_20_112 ();
 FILLCELL_X1 FILLER_0_20_116 ();
 FILLCELL_X4 FILLER_0_20_121 ();
 FILLCELL_X2 FILLER_0_20_125 ();
 FILLCELL_X1 FILLER_0_20_133 ();
 FILLCELL_X2 FILLER_0_20_163 ();
 FILLCELL_X8 FILLER_0_20_178 ();
 FILLCELL_X4 FILLER_0_20_186 ();
 FILLCELL_X4 FILLER_0_20_202 ();
 FILLCELL_X2 FILLER_0_20_206 ();
 FILLCELL_X1 FILLER_0_20_208 ();
 FILLCELL_X1 FILLER_0_20_225 ();
 FILLCELL_X4 FILLER_0_20_234 ();
 FILLCELL_X2 FILLER_0_20_238 ();
 FILLCELL_X2 FILLER_0_20_259 ();
 FILLCELL_X1 FILLER_0_20_261 ();
 FILLCELL_X2 FILLER_0_20_269 ();
 FILLCELL_X1 FILLER_0_20_278 ();
 FILLCELL_X2 FILLER_0_20_283 ();
 FILLCELL_X4 FILLER_0_20_290 ();
 FILLCELL_X2 FILLER_0_20_294 ();
 FILLCELL_X8 FILLER_0_20_307 ();
 FILLCELL_X4 FILLER_0_20_318 ();
 FILLCELL_X2 FILLER_0_20_322 ();
 FILLCELL_X1 FILLER_0_20_324 ();
 FILLCELL_X2 FILLER_0_20_333 ();
 FILLCELL_X1 FILLER_0_20_340 ();
 FILLCELL_X1 FILLER_0_20_354 ();
 FILLCELL_X1 FILLER_0_20_362 ();
 FILLCELL_X4 FILLER_0_20_372 ();
 FILLCELL_X1 FILLER_0_20_376 ();
 FILLCELL_X1 FILLER_0_20_380 ();
 FILLCELL_X4 FILLER_0_20_390 ();
 FILLCELL_X2 FILLER_0_20_408 ();
 FILLCELL_X1 FILLER_0_20_410 ();
 FILLCELL_X1 FILLER_0_21_16 ();
 FILLCELL_X1 FILLER_0_21_24 ();
 FILLCELL_X2 FILLER_0_21_27 ();
 FILLCELL_X2 FILLER_0_21_36 ();
 FILLCELL_X8 FILLER_0_21_42 ();
 FILLCELL_X1 FILLER_0_21_50 ();
 FILLCELL_X4 FILLER_0_21_54 ();
 FILLCELL_X2 FILLER_0_21_58 ();
 FILLCELL_X1 FILLER_0_21_60 ();
 FILLCELL_X2 FILLER_0_21_63 ();
 FILLCELL_X1 FILLER_0_21_65 ();
 FILLCELL_X2 FILLER_0_21_73 ();
 FILLCELL_X8 FILLER_0_21_77 ();
 FILLCELL_X1 FILLER_0_21_85 ();
 FILLCELL_X4 FILLER_0_21_90 ();
 FILLCELL_X2 FILLER_0_21_94 ();
 FILLCELL_X8 FILLER_0_21_113 ();
 FILLCELL_X4 FILLER_0_21_124 ();
 FILLCELL_X2 FILLER_0_21_128 ();
 FILLCELL_X2 FILLER_0_21_158 ();
 FILLCELL_X2 FILLER_0_21_223 ();
 FILLCELL_X8 FILLER_0_21_231 ();
 FILLCELL_X4 FILLER_0_21_239 ();
 FILLCELL_X2 FILLER_0_21_243 ();
 FILLCELL_X1 FILLER_0_21_245 ();
 FILLCELL_X1 FILLER_0_21_254 ();
 FILLCELL_X1 FILLER_0_21_259 ();
 FILLCELL_X4 FILLER_0_21_288 ();
 FILLCELL_X1 FILLER_0_21_302 ();
 FILLCELL_X2 FILLER_0_21_308 ();
 FILLCELL_X2 FILLER_0_21_315 ();
 FILLCELL_X2 FILLER_0_21_321 ();
 FILLCELL_X1 FILLER_0_21_323 ();
 FILLCELL_X1 FILLER_0_21_331 ();
 FILLCELL_X2 FILLER_0_21_345 ();
 FILLCELL_X4 FILLER_0_21_377 ();
 FILLCELL_X1 FILLER_0_21_381 ();
 FILLCELL_X4 FILLER_0_21_389 ();
 FILLCELL_X1 FILLER_0_21_393 ();
 FILLCELL_X2 FILLER_0_21_401 ();
 FILLCELL_X1 FILLER_0_21_403 ();
 FILLCELL_X1 FILLER_0_22_4 ();
 FILLCELL_X1 FILLER_0_22_8 ();
 FILLCELL_X1 FILLER_0_22_49 ();
 FILLCELL_X4 FILLER_0_22_54 ();
 FILLCELL_X2 FILLER_0_22_58 ();
 FILLCELL_X1 FILLER_0_22_60 ();
 FILLCELL_X4 FILLER_0_22_77 ();
 FILLCELL_X2 FILLER_0_22_93 ();
 FILLCELL_X1 FILLER_0_22_99 ();
 FILLCELL_X1 FILLER_0_22_140 ();
 FILLCELL_X8 FILLER_0_22_150 ();
 FILLCELL_X2 FILLER_0_22_158 ();
 FILLCELL_X1 FILLER_0_22_162 ();
 FILLCELL_X1 FILLER_0_22_166 ();
 FILLCELL_X1 FILLER_0_22_171 ();
 FILLCELL_X16 FILLER_0_22_176 ();
 FILLCELL_X8 FILLER_0_22_192 ();
 FILLCELL_X2 FILLER_0_22_208 ();
 FILLCELL_X8 FILLER_0_22_220 ();
 FILLCELL_X4 FILLER_0_22_228 ();
 FILLCELL_X2 FILLER_0_22_232 ();
 FILLCELL_X4 FILLER_0_22_238 ();
 FILLCELL_X1 FILLER_0_22_267 ();
 FILLCELL_X4 FILLER_0_22_293 ();
 FILLCELL_X2 FILLER_0_22_297 ();
 FILLCELL_X1 FILLER_0_22_299 ();
 FILLCELL_X1 FILLER_0_22_311 ();
 FILLCELL_X8 FILLER_0_22_317 ();
 FILLCELL_X2 FILLER_0_22_329 ();
 FILLCELL_X1 FILLER_0_22_331 ();
 FILLCELL_X4 FILLER_0_22_372 ();
 FILLCELL_X2 FILLER_0_22_376 ();
 FILLCELL_X2 FILLER_0_22_388 ();
 FILLCELL_X4 FILLER_0_22_396 ();
 FILLCELL_X4 FILLER_0_22_407 ();
 FILLCELL_X2 FILLER_0_23_1 ();
 FILLCELL_X8 FILLER_0_23_29 ();
 FILLCELL_X4 FILLER_0_23_37 ();
 FILLCELL_X2 FILLER_0_23_48 ();
 FILLCELL_X8 FILLER_0_23_66 ();
 FILLCELL_X2 FILLER_0_23_81 ();
 FILLCELL_X1 FILLER_0_23_83 ();
 FILLCELL_X1 FILLER_0_23_110 ();
 FILLCELL_X2 FILLER_0_23_116 ();
 FILLCELL_X1 FILLER_0_23_125 ();
 FILLCELL_X2 FILLER_0_23_129 ();
 FILLCELL_X8 FILLER_0_23_161 ();
 FILLCELL_X2 FILLER_0_23_169 ();
 FILLCELL_X16 FILLER_0_23_182 ();
 FILLCELL_X8 FILLER_0_23_198 ();
 FILLCELL_X1 FILLER_0_23_206 ();
 FILLCELL_X1 FILLER_0_23_214 ();
 FILLCELL_X8 FILLER_0_23_219 ();
 FILLCELL_X2 FILLER_0_23_227 ();
 FILLCELL_X2 FILLER_0_23_258 ();
 FILLCELL_X2 FILLER_0_23_267 ();
 FILLCELL_X1 FILLER_0_23_269 ();
 FILLCELL_X2 FILLER_0_23_273 ();
 FILLCELL_X1 FILLER_0_23_275 ();
 FILLCELL_X8 FILLER_0_23_287 ();
 FILLCELL_X8 FILLER_0_23_310 ();
 FILLCELL_X4 FILLER_0_23_341 ();
 FILLCELL_X4 FILLER_0_23_371 ();
 FILLCELL_X2 FILLER_0_23_375 ();
 FILLCELL_X1 FILLER_0_23_377 ();
 FILLCELL_X2 FILLER_0_23_394 ();
 FILLCELL_X1 FILLER_0_23_396 ();
 FILLCELL_X1 FILLER_0_24_4 ();
 FILLCELL_X1 FILLER_0_24_25 ();
 FILLCELL_X1 FILLER_0_24_30 ();
 FILLCELL_X8 FILLER_0_24_34 ();
 FILLCELL_X1 FILLER_0_24_42 ();
 FILLCELL_X4 FILLER_0_24_57 ();
 FILLCELL_X1 FILLER_0_24_61 ();
 FILLCELL_X4 FILLER_0_24_89 ();
 FILLCELL_X2 FILLER_0_24_98 ();
 FILLCELL_X1 FILLER_0_24_110 ();
 FILLCELL_X2 FILLER_0_24_119 ();
 FILLCELL_X2 FILLER_0_24_144 ();
 FILLCELL_X2 FILLER_0_24_155 ();
 FILLCELL_X1 FILLER_0_24_157 ();
 FILLCELL_X8 FILLER_0_24_188 ();
 FILLCELL_X2 FILLER_0_24_196 ();
 FILLCELL_X2 FILLER_0_24_207 ();
 FILLCELL_X2 FILLER_0_24_213 ();
 FILLCELL_X1 FILLER_0_24_215 ();
 FILLCELL_X4 FILLER_0_24_218 ();
 FILLCELL_X1 FILLER_0_24_222 ();
 FILLCELL_X2 FILLER_0_24_244 ();
 FILLCELL_X4 FILLER_0_24_253 ();
 FILLCELL_X2 FILLER_0_24_271 ();
 FILLCELL_X4 FILLER_0_24_280 ();
 FILLCELL_X2 FILLER_0_24_284 ();
 FILLCELL_X1 FILLER_0_24_286 ();
 FILLCELL_X1 FILLER_0_24_306 ();
 FILLCELL_X8 FILLER_0_24_313 ();
 FILLCELL_X1 FILLER_0_24_328 ();
 FILLCELL_X2 FILLER_0_24_336 ();
 FILLCELL_X4 FILLER_0_24_342 ();
 FILLCELL_X2 FILLER_0_24_373 ();
 FILLCELL_X1 FILLER_0_24_375 ();
 FILLCELL_X2 FILLER_0_24_383 ();
 FILLCELL_X2 FILLER_0_24_389 ();
 FILLCELL_X1 FILLER_0_24_391 ();
 FILLCELL_X4 FILLER_0_24_406 ();
 FILLCELL_X1 FILLER_0_24_410 ();
 FILLCELL_X1 FILLER_0_25_7 ();
 FILLCELL_X2 FILLER_0_25_16 ();
 FILLCELL_X1 FILLER_0_25_18 ();
 FILLCELL_X2 FILLER_0_25_23 ();
 FILLCELL_X1 FILLER_0_25_25 ();
 FILLCELL_X4 FILLER_0_25_29 ();
 FILLCELL_X1 FILLER_0_25_33 ();
 FILLCELL_X1 FILLER_0_25_42 ();
 FILLCELL_X1 FILLER_0_25_53 ();
 FILLCELL_X1 FILLER_0_25_61 ();
 FILLCELL_X1 FILLER_0_25_65 ();
 FILLCELL_X2 FILLER_0_25_75 ();
 FILLCELL_X2 FILLER_0_25_80 ();
 FILLCELL_X1 FILLER_0_25_96 ();
 FILLCELL_X1 FILLER_0_25_101 ();
 FILLCELL_X1 FILLER_0_25_111 ();
 FILLCELL_X2 FILLER_0_25_117 ();
 FILLCELL_X2 FILLER_0_25_122 ();
 FILLCELL_X2 FILLER_0_25_146 ();
 FILLCELL_X4 FILLER_0_25_158 ();
 FILLCELL_X16 FILLER_0_25_187 ();
 FILLCELL_X4 FILLER_0_25_203 ();
 FILLCELL_X2 FILLER_0_25_207 ();
 FILLCELL_X1 FILLER_0_25_209 ();
 FILLCELL_X8 FILLER_0_25_219 ();
 FILLCELL_X4 FILLER_0_25_227 ();
 FILLCELL_X2 FILLER_0_25_231 ();
 FILLCELL_X8 FILLER_0_25_240 ();
 FILLCELL_X4 FILLER_0_25_248 ();
 FILLCELL_X1 FILLER_0_25_252 ();
 FILLCELL_X2 FILLER_0_25_260 ();
 FILLCELL_X1 FILLER_0_25_262 ();
 FILLCELL_X2 FILLER_0_25_277 ();
 FILLCELL_X8 FILLER_0_25_284 ();
 FILLCELL_X4 FILLER_0_25_292 ();
 FILLCELL_X2 FILLER_0_25_296 ();
 FILLCELL_X1 FILLER_0_25_298 ();
 FILLCELL_X8 FILLER_0_25_308 ();
 FILLCELL_X2 FILLER_0_25_316 ();
 FILLCELL_X1 FILLER_0_25_318 ();
 FILLCELL_X4 FILLER_0_25_332 ();
 FILLCELL_X1 FILLER_0_25_336 ();
 FILLCELL_X1 FILLER_0_25_379 ();
 FILLCELL_X1 FILLER_0_25_396 ();
 FILLCELL_X4 FILLER_0_26_1 ();
 FILLCELL_X1 FILLER_0_26_5 ();
 FILLCELL_X1 FILLER_0_26_13 ();
 FILLCELL_X2 FILLER_0_26_25 ();
 FILLCELL_X1 FILLER_0_26_30 ();
 FILLCELL_X4 FILLER_0_26_41 ();
 FILLCELL_X4 FILLER_0_26_49 ();
 FILLCELL_X1 FILLER_0_26_53 ();
 FILLCELL_X4 FILLER_0_26_80 ();
 FILLCELL_X1 FILLER_0_26_84 ();
 FILLCELL_X8 FILLER_0_26_94 ();
 FILLCELL_X1 FILLER_0_26_106 ();
 FILLCELL_X1 FILLER_0_26_111 ();
 FILLCELL_X1 FILLER_0_26_119 ();
 FILLCELL_X1 FILLER_0_26_150 ();
 FILLCELL_X2 FILLER_0_26_157 ();
 FILLCELL_X1 FILLER_0_26_159 ();
 FILLCELL_X1 FILLER_0_26_170 ();
 FILLCELL_X1 FILLER_0_26_176 ();
 FILLCELL_X1 FILLER_0_26_182 ();
 FILLCELL_X2 FILLER_0_26_187 ();
 FILLCELL_X1 FILLER_0_26_189 ();
 FILLCELL_X4 FILLER_0_26_209 ();
 FILLCELL_X4 FILLER_0_26_218 ();
 FILLCELL_X1 FILLER_0_26_222 ();
 FILLCELL_X4 FILLER_0_26_235 ();
 FILLCELL_X1 FILLER_0_26_243 ();
 FILLCELL_X4 FILLER_0_26_258 ();
 FILLCELL_X1 FILLER_0_26_262 ();
 FILLCELL_X8 FILLER_0_26_287 ();
 FILLCELL_X4 FILLER_0_26_295 ();
 FILLCELL_X2 FILLER_0_26_299 ();
 FILLCELL_X1 FILLER_0_26_301 ();
 FILLCELL_X8 FILLER_0_26_307 ();
 FILLCELL_X1 FILLER_0_26_315 ();
 FILLCELL_X2 FILLER_0_26_340 ();
 FILLCELL_X2 FILLER_0_26_352 ();
 FILLCELL_X1 FILLER_0_26_357 ();
 FILLCELL_X2 FILLER_0_26_378 ();
 FILLCELL_X1 FILLER_0_26_403 ();
 FILLCELL_X8 FILLER_0_27_1 ();
 FILLCELL_X4 FILLER_0_27_9 ();
 FILLCELL_X1 FILLER_0_27_20 ();
 FILLCELL_X2 FILLER_0_27_39 ();
 FILLCELL_X1 FILLER_0_27_41 ();
 FILLCELL_X4 FILLER_0_27_49 ();
 FILLCELL_X2 FILLER_0_27_57 ();
 FILLCELL_X4 FILLER_0_27_65 ();
 FILLCELL_X1 FILLER_0_27_69 ();
 FILLCELL_X1 FILLER_0_27_95 ();
 FILLCELL_X4 FILLER_0_27_113 ();
 FILLCELL_X2 FILLER_0_27_219 ();
 FILLCELL_X2 FILLER_0_27_223 ();
 FILLCELL_X8 FILLER_0_27_232 ();
 FILLCELL_X1 FILLER_0_27_243 ();
 FILLCELL_X2 FILLER_0_27_248 ();
 FILLCELL_X1 FILLER_0_27_250 ();
 FILLCELL_X4 FILLER_0_27_258 ();
 FILLCELL_X1 FILLER_0_27_262 ();
 FILLCELL_X1 FILLER_0_27_270 ();
 FILLCELL_X2 FILLER_0_27_276 ();
 FILLCELL_X1 FILLER_0_27_278 ();
 FILLCELL_X8 FILLER_0_27_283 ();
 FILLCELL_X4 FILLER_0_27_291 ();
 FILLCELL_X2 FILLER_0_27_295 ();
 FILLCELL_X2 FILLER_0_27_302 ();
 FILLCELL_X1 FILLER_0_27_304 ();
 FILLCELL_X1 FILLER_0_27_310 ();
 FILLCELL_X2 FILLER_0_27_343 ();
 FILLCELL_X1 FILLER_0_27_345 ();
 FILLCELL_X1 FILLER_0_27_356 ();
 FILLCELL_X2 FILLER_0_27_360 ();
 FILLCELL_X2 FILLER_0_27_380 ();
 FILLCELL_X1 FILLER_0_27_386 ();
 FILLCELL_X2 FILLER_0_27_390 ();
 FILLCELL_X4 FILLER_0_27_399 ();
 FILLCELL_X1 FILLER_0_27_403 ();
 FILLCELL_X8 FILLER_0_28_1 ();
 FILLCELL_X4 FILLER_0_28_9 ();
 FILLCELL_X2 FILLER_0_28_22 ();
 FILLCELL_X2 FILLER_0_28_31 ();
 FILLCELL_X2 FILLER_0_28_37 ();
 FILLCELL_X8 FILLER_0_28_48 ();
 FILLCELL_X2 FILLER_0_28_62 ();
 FILLCELL_X1 FILLER_0_28_64 ();
 FILLCELL_X8 FILLER_0_28_71 ();
 FILLCELL_X1 FILLER_0_28_79 ();
 FILLCELL_X2 FILLER_0_28_95 ();
 FILLCELL_X1 FILLER_0_28_104 ();
 FILLCELL_X1 FILLER_0_28_116 ();
 FILLCELL_X8 FILLER_0_28_127 ();
 FILLCELL_X4 FILLER_0_28_135 ();
 FILLCELL_X1 FILLER_0_28_146 ();
 FILLCELL_X2 FILLER_0_28_156 ();
 FILLCELL_X4 FILLER_0_28_162 ();
 FILLCELL_X32 FILLER_0_28_168 ();
 FILLCELL_X4 FILLER_0_28_200 ();
 FILLCELL_X1 FILLER_0_28_204 ();
 FILLCELL_X8 FILLER_0_28_215 ();
 FILLCELL_X2 FILLER_0_28_223 ();
 FILLCELL_X4 FILLER_0_28_232 ();
 FILLCELL_X2 FILLER_0_28_236 ();
 FILLCELL_X1 FILLER_0_28_259 ();
 FILLCELL_X2 FILLER_0_28_282 ();
 FILLCELL_X4 FILLER_0_28_294 ();
 FILLCELL_X2 FILLER_0_28_314 ();
 FILLCELL_X2 FILLER_0_28_347 ();
 FILLCELL_X2 FILLER_0_28_353 ();
 FILLCELL_X2 FILLER_0_28_360 ();
 FILLCELL_X1 FILLER_0_28_362 ();
 FILLCELL_X4 FILLER_0_28_399 ();
 FILLCELL_X1 FILLER_0_28_403 ();
 FILLCELL_X2 FILLER_0_29_1 ();
 FILLCELL_X1 FILLER_0_29_3 ();
 FILLCELL_X1 FILLER_0_29_22 ();
 FILLCELL_X1 FILLER_0_29_27 ();
 FILLCELL_X1 FILLER_0_29_32 ();
 FILLCELL_X2 FILLER_0_29_36 ();
 FILLCELL_X1 FILLER_0_29_47 ();
 FILLCELL_X1 FILLER_0_29_52 ();
 FILLCELL_X4 FILLER_0_29_79 ();
 FILLCELL_X2 FILLER_0_29_83 ();
 FILLCELL_X1 FILLER_0_29_85 ();
 FILLCELL_X2 FILLER_0_29_109 ();
 FILLCELL_X2 FILLER_0_29_114 ();
 FILLCELL_X2 FILLER_0_29_132 ();
 FILLCELL_X1 FILLER_0_29_134 ();
 FILLCELL_X2 FILLER_0_29_138 ();
 FILLCELL_X1 FILLER_0_29_140 ();
 FILLCELL_X8 FILLER_0_29_156 ();
 FILLCELL_X1 FILLER_0_29_164 ();
 FILLCELL_X1 FILLER_0_29_174 ();
 FILLCELL_X2 FILLER_0_29_191 ();
 FILLCELL_X1 FILLER_0_29_193 ();
 FILLCELL_X2 FILLER_0_29_209 ();
 FILLCELL_X1 FILLER_0_29_226 ();
 FILLCELL_X4 FILLER_0_29_259 ();
 FILLCELL_X2 FILLER_0_29_263 ();
 FILLCELL_X1 FILLER_0_29_279 ();
 FILLCELL_X4 FILLER_0_29_284 ();
 FILLCELL_X16 FILLER_0_29_303 ();
 FILLCELL_X4 FILLER_0_29_319 ();
 FILLCELL_X2 FILLER_0_29_323 ();
 FILLCELL_X4 FILLER_0_29_395 ();
 FILLCELL_X4 FILLER_0_29_406 ();
 FILLCELL_X1 FILLER_0_29_410 ();
 FILLCELL_X8 FILLER_0_30_1 ();
 FILLCELL_X1 FILLER_0_30_9 ();
 FILLCELL_X1 FILLER_0_30_18 ();
 FILLCELL_X4 FILLER_0_30_34 ();
 FILLCELL_X1 FILLER_0_30_38 ();
 FILLCELL_X2 FILLER_0_30_43 ();
 FILLCELL_X4 FILLER_0_30_49 ();
 FILLCELL_X2 FILLER_0_30_53 ();
 FILLCELL_X2 FILLER_0_30_59 ();
 FILLCELL_X1 FILLER_0_30_61 ();
 FILLCELL_X8 FILLER_0_30_66 ();
 FILLCELL_X2 FILLER_0_30_74 ();
 FILLCELL_X4 FILLER_0_30_80 ();
 FILLCELL_X1 FILLER_0_30_84 ();
 FILLCELL_X2 FILLER_0_30_88 ();
 FILLCELL_X1 FILLER_0_30_90 ();
 FILLCELL_X8 FILLER_0_30_152 ();
 FILLCELL_X4 FILLER_0_30_160 ();
 FILLCELL_X2 FILLER_0_30_164 ();
 FILLCELL_X1 FILLER_0_30_186 ();
 FILLCELL_X16 FILLER_0_30_192 ();
 FILLCELL_X2 FILLER_0_30_215 ();
 FILLCELL_X4 FILLER_0_30_220 ();
 FILLCELL_X8 FILLER_0_30_253 ();
 FILLCELL_X1 FILLER_0_30_261 ();
 FILLCELL_X8 FILLER_0_30_282 ();
 FILLCELL_X4 FILLER_0_30_290 ();
 FILLCELL_X8 FILLER_0_30_305 ();
 FILLCELL_X2 FILLER_0_30_313 ();
 FILLCELL_X1 FILLER_0_30_321 ();
 FILLCELL_X2 FILLER_0_30_325 ();
 FILLCELL_X1 FILLER_0_30_327 ();
 FILLCELL_X1 FILLER_0_30_332 ();
 FILLCELL_X2 FILLER_0_30_358 ();
 FILLCELL_X2 FILLER_0_30_364 ();
 FILLCELL_X2 FILLER_0_30_374 ();
 FILLCELL_X1 FILLER_0_30_383 ();
 FILLCELL_X1 FILLER_0_30_387 ();
 FILLCELL_X1 FILLER_0_30_394 ();
 FILLCELL_X2 FILLER_0_30_402 ();
 FILLCELL_X8 FILLER_0_31_1 ();
 FILLCELL_X4 FILLER_0_31_9 ();
 FILLCELL_X1 FILLER_0_31_13 ();
 FILLCELL_X4 FILLER_0_31_21 ();
 FILLCELL_X1 FILLER_0_31_25 ();
 FILLCELL_X2 FILLER_0_31_32 ();
 FILLCELL_X1 FILLER_0_31_34 ();
 FILLCELL_X1 FILLER_0_31_37 ();
 FILLCELL_X2 FILLER_0_31_41 ();
 FILLCELL_X2 FILLER_0_31_67 ();
 FILLCELL_X8 FILLER_0_31_73 ();
 FILLCELL_X1 FILLER_0_31_81 ();
 FILLCELL_X1 FILLER_0_31_86 ();
 FILLCELL_X1 FILLER_0_31_89 ();
 FILLCELL_X1 FILLER_0_31_94 ();
 FILLCELL_X1 FILLER_0_31_106 ();
 FILLCELL_X1 FILLER_0_31_109 ();
 FILLCELL_X4 FILLER_0_31_121 ();
 FILLCELL_X2 FILLER_0_31_125 ();
 FILLCELL_X1 FILLER_0_31_127 ();
 FILLCELL_X1 FILLER_0_31_158 ();
 FILLCELL_X1 FILLER_0_31_165 ();
 FILLCELL_X1 FILLER_0_31_176 ();
 FILLCELL_X1 FILLER_0_31_185 ();
 FILLCELL_X16 FILLER_0_31_190 ();
 FILLCELL_X4 FILLER_0_31_206 ();
 FILLCELL_X2 FILLER_0_31_210 ();
 FILLCELL_X16 FILLER_0_31_223 ();
 FILLCELL_X8 FILLER_0_31_260 ();
 FILLCELL_X2 FILLER_0_31_268 ();
 FILLCELL_X1 FILLER_0_31_270 ();
 FILLCELL_X8 FILLER_0_31_280 ();
 FILLCELL_X4 FILLER_0_31_288 ();
 FILLCELL_X1 FILLER_0_31_319 ();
 FILLCELL_X4 FILLER_0_31_324 ();
 FILLCELL_X2 FILLER_0_31_328 ();
 FILLCELL_X4 FILLER_0_31_345 ();
 FILLCELL_X1 FILLER_0_31_349 ();
 FILLCELL_X8 FILLER_0_31_362 ();
 FILLCELL_X4 FILLER_0_31_370 ();
 FILLCELL_X2 FILLER_0_31_374 ();
 FILLCELL_X2 FILLER_0_31_379 ();
 FILLCELL_X1 FILLER_0_31_391 ();
 FILLCELL_X4 FILLER_0_31_399 ();
 FILLCELL_X1 FILLER_0_31_403 ();
 FILLCELL_X2 FILLER_0_32_1 ();
 FILLCELL_X1 FILLER_0_32_3 ();
 FILLCELL_X1 FILLER_0_32_6 ();
 FILLCELL_X1 FILLER_0_32_11 ();
 FILLCELL_X1 FILLER_0_32_19 ();
 FILLCELL_X1 FILLER_0_32_30 ();
 FILLCELL_X1 FILLER_0_32_35 ();
 FILLCELL_X1 FILLER_0_32_41 ();
 FILLCELL_X1 FILLER_0_32_47 ();
 FILLCELL_X1 FILLER_0_32_54 ();
 FILLCELL_X2 FILLER_0_32_60 ();
 FILLCELL_X8 FILLER_0_32_66 ();
 FILLCELL_X4 FILLER_0_32_74 ();
 FILLCELL_X2 FILLER_0_32_78 ();
 FILLCELL_X1 FILLER_0_32_80 ();
 FILLCELL_X2 FILLER_0_32_148 ();
 FILLCELL_X4 FILLER_0_32_154 ();
 FILLCELL_X2 FILLER_0_32_158 ();
 FILLCELL_X2 FILLER_0_32_198 ();
 FILLCELL_X1 FILLER_0_32_200 ();
 FILLCELL_X1 FILLER_0_32_223 ();
 FILLCELL_X2 FILLER_0_32_227 ();
 FILLCELL_X4 FILLER_0_32_261 ();
 FILLCELL_X2 FILLER_0_32_265 ();
 FILLCELL_X2 FILLER_0_32_301 ();
 FILLCELL_X1 FILLER_0_32_303 ();
 FILLCELL_X1 FILLER_0_32_309 ();
 FILLCELL_X1 FILLER_0_32_317 ();
 FILLCELL_X4 FILLER_0_32_325 ();
 FILLCELL_X1 FILLER_0_32_329 ();
 FILLCELL_X2 FILLER_0_32_337 ();
 FILLCELL_X8 FILLER_0_32_392 ();
 FILLCELL_X4 FILLER_0_32_400 ();
 FILLCELL_X16 FILLER_0_33_1 ();
 FILLCELL_X1 FILLER_0_33_25 ();
 FILLCELL_X1 FILLER_0_33_41 ();
 FILLCELL_X1 FILLER_0_33_51 ();
 FILLCELL_X1 FILLER_0_33_56 ();
 FILLCELL_X1 FILLER_0_33_91 ();
 FILLCELL_X2 FILLER_0_33_140 ();
 FILLCELL_X2 FILLER_0_33_145 ();
 FILLCELL_X2 FILLER_0_33_169 ();
 FILLCELL_X32 FILLER_0_33_179 ();
 FILLCELL_X1 FILLER_0_33_211 ();
 FILLCELL_X2 FILLER_0_33_215 ();
 FILLCELL_X2 FILLER_0_33_226 ();
 FILLCELL_X1 FILLER_0_33_228 ();
 FILLCELL_X2 FILLER_0_33_239 ();
 FILLCELL_X2 FILLER_0_33_245 ();
 FILLCELL_X1 FILLER_0_33_247 ();
 FILLCELL_X8 FILLER_0_33_255 ();
 FILLCELL_X1 FILLER_0_33_274 ();
 FILLCELL_X2 FILLER_0_33_292 ();
 FILLCELL_X1 FILLER_0_33_294 ();
 FILLCELL_X4 FILLER_0_33_299 ();
 FILLCELL_X2 FILLER_0_33_332 ();
 FILLCELL_X1 FILLER_0_33_370 ();
 FILLCELL_X2 FILLER_0_33_397 ();
 FILLCELL_X4 FILLER_0_33_406 ();
 FILLCELL_X1 FILLER_0_33_410 ();
 FILLCELL_X2 FILLER_0_34_5 ();
 FILLCELL_X1 FILLER_0_34_14 ();
 FILLCELL_X4 FILLER_0_34_24 ();
 FILLCELL_X2 FILLER_0_34_33 ();
 FILLCELL_X1 FILLER_0_34_46 ();
 FILLCELL_X2 FILLER_0_34_63 ();
 FILLCELL_X4 FILLER_0_34_71 ();
 FILLCELL_X2 FILLER_0_34_75 ();
 FILLCELL_X1 FILLER_0_34_87 ();
 FILLCELL_X4 FILLER_0_34_101 ();
 FILLCELL_X2 FILLER_0_34_152 ();
 FILLCELL_X16 FILLER_0_34_178 ();
 FILLCELL_X8 FILLER_0_34_194 ();
 FILLCELL_X4 FILLER_0_34_202 ();
 FILLCELL_X2 FILLER_0_34_206 ();
 FILLCELL_X1 FILLER_0_34_208 ();
 FILLCELL_X8 FILLER_0_34_229 ();
 FILLCELL_X2 FILLER_0_34_237 ();
 FILLCELL_X4 FILLER_0_34_248 ();
 FILLCELL_X2 FILLER_0_34_252 ();
 FILLCELL_X1 FILLER_0_34_254 ();
 FILLCELL_X1 FILLER_0_34_266 ();
 FILLCELL_X4 FILLER_0_34_274 ();
 FILLCELL_X2 FILLER_0_34_287 ();
 FILLCELL_X1 FILLER_0_34_314 ();
 FILLCELL_X8 FILLER_0_34_325 ();
 FILLCELL_X2 FILLER_0_34_347 ();
 FILLCELL_X2 FILLER_0_34_359 ();
 FILLCELL_X1 FILLER_0_34_361 ();
 FILLCELL_X4 FILLER_0_34_369 ();
 FILLCELL_X1 FILLER_0_34_373 ();
 FILLCELL_X1 FILLER_0_34_378 ();
 FILLCELL_X4 FILLER_0_34_399 ();
 FILLCELL_X1 FILLER_0_34_403 ();
 FILLCELL_X2 FILLER_0_35_1 ();
 FILLCELL_X1 FILLER_0_35_3 ();
 FILLCELL_X32 FILLER_0_35_33 ();
 FILLCELL_X8 FILLER_0_35_65 ();
 FILLCELL_X2 FILLER_0_35_73 ();
 FILLCELL_X4 FILLER_0_35_82 ();
 FILLCELL_X8 FILLER_0_35_99 ();
 FILLCELL_X2 FILLER_0_35_107 ();
 FILLCELL_X1 FILLER_0_35_118 ();
 FILLCELL_X1 FILLER_0_35_125 ();
 FILLCELL_X16 FILLER_0_35_133 ();
 FILLCELL_X4 FILLER_0_35_149 ();
 FILLCELL_X1 FILLER_0_35_153 ();
 FILLCELL_X2 FILLER_0_35_166 ();
 FILLCELL_X1 FILLER_0_35_168 ();
 FILLCELL_X4 FILLER_0_35_173 ();
 FILLCELL_X1 FILLER_0_35_177 ();
 FILLCELL_X4 FILLER_0_35_181 ();
 FILLCELL_X8 FILLER_0_35_201 ();
 FILLCELL_X1 FILLER_0_35_209 ();
 FILLCELL_X4 FILLER_0_35_221 ();
 FILLCELL_X4 FILLER_0_35_229 ();
 FILLCELL_X1 FILLER_0_35_233 ();
 FILLCELL_X1 FILLER_0_35_247 ();
 FILLCELL_X4 FILLER_0_35_291 ();
 FILLCELL_X2 FILLER_0_35_324 ();
 FILLCELL_X4 FILLER_0_35_341 ();
 FILLCELL_X4 FILLER_0_35_349 ();
 FILLCELL_X2 FILLER_0_35_353 ();
 FILLCELL_X4 FILLER_0_35_383 ();
 FILLCELL_X2 FILLER_0_35_387 ();
 FILLCELL_X1 FILLER_0_35_389 ();
 FILLCELL_X2 FILLER_0_36_28 ();
 FILLCELL_X1 FILLER_0_36_33 ();
 FILLCELL_X16 FILLER_0_36_38 ();
 FILLCELL_X4 FILLER_0_36_54 ();
 FILLCELL_X2 FILLER_0_36_58 ();
 FILLCELL_X1 FILLER_0_36_60 ();
 FILLCELL_X4 FILLER_0_36_99 ();
 FILLCELL_X1 FILLER_0_36_103 ();
 FILLCELL_X1 FILLER_0_36_112 ();
 FILLCELL_X2 FILLER_0_36_117 ();
 FILLCELL_X1 FILLER_0_36_119 ();
 FILLCELL_X16 FILLER_0_36_124 ();
 FILLCELL_X4 FILLER_0_36_156 ();
 FILLCELL_X2 FILLER_0_36_160 ();
 FILLCELL_X1 FILLER_0_36_162 ();
 FILLCELL_X1 FILLER_0_36_167 ();
 FILLCELL_X1 FILLER_0_36_207 ();
 FILLCELL_X1 FILLER_0_36_237 ();
 FILLCELL_X1 FILLER_0_36_243 ();
 FILLCELL_X2 FILLER_0_36_263 ();
 FILLCELL_X2 FILLER_0_36_292 ();
 FILLCELL_X2 FILLER_0_36_297 ();
 FILLCELL_X1 FILLER_0_36_307 ();
 FILLCELL_X1 FILLER_0_36_312 ();
 FILLCELL_X1 FILLER_0_36_321 ();
 FILLCELL_X32 FILLER_0_36_326 ();
 FILLCELL_X2 FILLER_0_36_358 ();
 FILLCELL_X1 FILLER_0_36_360 ();
 FILLCELL_X2 FILLER_0_36_363 ();
 FILLCELL_X1 FILLER_0_36_374 ();
 FILLCELL_X1 FILLER_0_36_392 ();
 FILLCELL_X4 FILLER_0_36_406 ();
 FILLCELL_X1 FILLER_0_36_410 ();
 FILLCELL_X1 FILLER_0_37_8 ();
 FILLCELL_X1 FILLER_0_37_17 ();
 FILLCELL_X1 FILLER_0_37_22 ();
 FILLCELL_X1 FILLER_0_37_30 ();
 FILLCELL_X2 FILLER_0_37_34 ();
 FILLCELL_X1 FILLER_0_37_53 ();
 FILLCELL_X2 FILLER_0_37_88 ();
 FILLCELL_X4 FILLER_0_37_96 ();
 FILLCELL_X2 FILLER_0_37_100 ();
 FILLCELL_X2 FILLER_0_37_109 ();
 FILLCELL_X4 FILLER_0_37_117 ();
 FILLCELL_X2 FILLER_0_37_121 ();
 FILLCELL_X1 FILLER_0_37_123 ();
 FILLCELL_X8 FILLER_0_37_183 ();
 FILLCELL_X4 FILLER_0_37_191 ();
 FILLCELL_X2 FILLER_0_37_204 ();
 FILLCELL_X4 FILLER_0_37_233 ();
 FILLCELL_X1 FILLER_0_37_237 ();
 FILLCELL_X8 FILLER_0_37_245 ();
 FILLCELL_X2 FILLER_0_37_253 ();
 FILLCELL_X1 FILLER_0_37_269 ();
 FILLCELL_X4 FILLER_0_37_295 ();
 FILLCELL_X1 FILLER_0_37_299 ();
 FILLCELL_X2 FILLER_0_37_311 ();
 FILLCELL_X32 FILLER_0_37_317 ();
 FILLCELL_X8 FILLER_0_37_349 ();
 FILLCELL_X4 FILLER_0_37_357 ();
 FILLCELL_X1 FILLER_0_37_377 ();
 FILLCELL_X2 FILLER_0_37_385 ();
 FILLCELL_X1 FILLER_0_37_394 ();
 FILLCELL_X2 FILLER_0_37_402 ();
 FILLCELL_X2 FILLER_0_38_34 ();
 FILLCELL_X2 FILLER_0_38_40 ();
 FILLCELL_X1 FILLER_0_38_73 ();
 FILLCELL_X1 FILLER_0_38_78 ();
 FILLCELL_X1 FILLER_0_38_83 ();
 FILLCELL_X8 FILLER_0_38_112 ();
 FILLCELL_X4 FILLER_0_38_120 ();
 FILLCELL_X2 FILLER_0_38_124 ();
 FILLCELL_X4 FILLER_0_38_147 ();
 FILLCELL_X1 FILLER_0_38_161 ();
 FILLCELL_X1 FILLER_0_38_170 ();
 FILLCELL_X1 FILLER_0_38_173 ();
 FILLCELL_X1 FILLER_0_38_180 ();
 FILLCELL_X1 FILLER_0_38_197 ();
 FILLCELL_X4 FILLER_0_38_217 ();
 FILLCELL_X1 FILLER_0_38_226 ();
 FILLCELL_X2 FILLER_0_38_230 ();
 FILLCELL_X4 FILLER_0_38_236 ();
 FILLCELL_X32 FILLER_0_38_300 ();
 FILLCELL_X32 FILLER_0_38_332 ();
 FILLCELL_X8 FILLER_0_38_364 ();
 FILLCELL_X4 FILLER_0_38_372 ();
 FILLCELL_X1 FILLER_0_38_376 ();
 FILLCELL_X4 FILLER_0_38_398 ();
 FILLCELL_X2 FILLER_0_38_402 ();
 FILLCELL_X1 FILLER_0_39_13 ();
 FILLCELL_X1 FILLER_0_39_38 ();
 FILLCELL_X4 FILLER_0_39_46 ();
 FILLCELL_X1 FILLER_0_39_50 ();
 FILLCELL_X2 FILLER_0_39_77 ();
 FILLCELL_X1 FILLER_0_39_89 ();
 FILLCELL_X1 FILLER_0_39_112 ();
 FILLCELL_X4 FILLER_0_39_119 ();
 FILLCELL_X2 FILLER_0_39_123 ();
 FILLCELL_X8 FILLER_0_39_144 ();
 FILLCELL_X2 FILLER_0_39_152 ();
 FILLCELL_X1 FILLER_0_39_166 ();
 FILLCELL_X4 FILLER_0_39_187 ();
 FILLCELL_X8 FILLER_0_39_207 ();
 FILLCELL_X1 FILLER_0_39_215 ();
 FILLCELL_X2 FILLER_0_39_222 ();
 FILLCELL_X1 FILLER_0_39_224 ();
 FILLCELL_X1 FILLER_0_39_236 ();
 FILLCELL_X4 FILLER_0_39_244 ();
 FILLCELL_X2 FILLER_0_39_248 ();
 FILLCELL_X1 FILLER_0_39_250 ();
 FILLCELL_X4 FILLER_0_39_258 ();
 FILLCELL_X2 FILLER_0_39_262 ();
 FILLCELL_X32 FILLER_0_39_269 ();
 FILLCELL_X32 FILLER_0_39_301 ();
 FILLCELL_X32 FILLER_0_39_333 ();
 FILLCELL_X16 FILLER_0_39_365 ();
 FILLCELL_X8 FILLER_0_39_381 ();
 FILLCELL_X1 FILLER_0_39_389 ();
 FILLCELL_X1 FILLER_0_40_20 ();
 FILLCELL_X1 FILLER_0_40_56 ();
 FILLCELL_X2 FILLER_0_40_61 ();
 FILLCELL_X2 FILLER_0_40_74 ();
 FILLCELL_X1 FILLER_0_40_106 ();
 FILLCELL_X16 FILLER_0_40_113 ();
 FILLCELL_X4 FILLER_0_40_139 ();
 FILLCELL_X2 FILLER_0_40_143 ();
 FILLCELL_X1 FILLER_0_40_145 ();
 FILLCELL_X1 FILLER_0_40_148 ();
 FILLCELL_X2 FILLER_0_40_182 ();
 FILLCELL_X4 FILLER_0_40_186 ();
 FILLCELL_X1 FILLER_0_40_190 ();
 FILLCELL_X4 FILLER_0_40_207 ();
 FILLCELL_X2 FILLER_0_40_211 ();
 FILLCELL_X32 FILLER_0_40_223 ();
 FILLCELL_X32 FILLER_0_40_255 ();
 FILLCELL_X32 FILLER_0_40_287 ();
 FILLCELL_X32 FILLER_0_40_319 ();
 FILLCELL_X32 FILLER_0_40_351 ();
 FILLCELL_X16 FILLER_0_40_383 ();
 FILLCELL_X8 FILLER_0_40_399 ();
 FILLCELL_X4 FILLER_0_40_407 ();
 FILLCELL_X1 FILLER_0_41_1 ();
 FILLCELL_X1 FILLER_0_41_10 ();
 FILLCELL_X1 FILLER_0_41_19 ();
 FILLCELL_X2 FILLER_0_41_23 ();
 FILLCELL_X32 FILLER_0_41_28 ();
 FILLCELL_X32 FILLER_0_41_60 ();
 FILLCELL_X16 FILLER_0_41_92 ();
 FILLCELL_X2 FILLER_0_41_108 ();
 FILLCELL_X16 FILLER_0_41_120 ();
 FILLCELL_X4 FILLER_0_41_136 ();
 FILLCELL_X4 FILLER_0_41_150 ();
 FILLCELL_X4 FILLER_0_41_156 ();
 FILLCELL_X32 FILLER_0_41_196 ();
 FILLCELL_X32 FILLER_0_41_228 ();
 FILLCELL_X32 FILLER_0_41_260 ();
 FILLCELL_X32 FILLER_0_41_292 ();
 FILLCELL_X32 FILLER_0_41_324 ();
 FILLCELL_X32 FILLER_0_41_356 ();
 FILLCELL_X16 FILLER_0_41_388 ();
 FILLCELL_X4 FILLER_0_41_404 ();
 FILLCELL_X2 FILLER_0_41_408 ();
 FILLCELL_X1 FILLER_0_41_410 ();
 FILLCELL_X2 FILLER_0_42_1 ();
 FILLCELL_X32 FILLER_0_42_7 ();
 FILLCELL_X32 FILLER_0_42_39 ();
 FILLCELL_X32 FILLER_0_42_71 ();
 FILLCELL_X32 FILLER_0_42_103 ();
 FILLCELL_X16 FILLER_0_42_135 ();
 FILLCELL_X8 FILLER_0_42_151 ();
 FILLCELL_X4 FILLER_0_42_159 ();
 FILLCELL_X2 FILLER_0_42_163 ();
 FILLCELL_X1 FILLER_0_42_165 ();
 FILLCELL_X32 FILLER_0_42_168 ();
 FILLCELL_X32 FILLER_0_42_200 ();
 FILLCELL_X32 FILLER_0_42_232 ();
 FILLCELL_X32 FILLER_0_42_264 ();
 FILLCELL_X32 FILLER_0_42_296 ();
 FILLCELL_X32 FILLER_0_42_328 ();
 FILLCELL_X32 FILLER_0_42_360 ();
 FILLCELL_X16 FILLER_0_42_392 ();
 FILLCELL_X2 FILLER_0_42_408 ();
 FILLCELL_X1 FILLER_0_42_410 ();
 FILLCELL_X32 FILLER_0_43_1 ();
 FILLCELL_X32 FILLER_0_43_33 ();
 FILLCELL_X32 FILLER_0_43_65 ();
 FILLCELL_X32 FILLER_0_43_97 ();
 FILLCELL_X32 FILLER_0_43_129 ();
 FILLCELL_X32 FILLER_0_43_161 ();
 FILLCELL_X32 FILLER_0_43_193 ();
 FILLCELL_X32 FILLER_0_43_225 ();
 FILLCELL_X32 FILLER_0_43_257 ();
 FILLCELL_X32 FILLER_0_43_289 ();
 FILLCELL_X32 FILLER_0_43_321 ();
 FILLCELL_X32 FILLER_0_43_353 ();
 FILLCELL_X16 FILLER_0_43_385 ();
 FILLCELL_X8 FILLER_0_43_401 ();
 FILLCELL_X2 FILLER_0_43_409 ();
 FILLCELL_X32 FILLER_0_44_1 ();
 FILLCELL_X32 FILLER_0_44_33 ();
 FILLCELL_X32 FILLER_0_44_65 ();
 FILLCELL_X32 FILLER_0_44_97 ();
 FILLCELL_X32 FILLER_0_44_129 ();
 FILLCELL_X32 FILLER_0_44_161 ();
 FILLCELL_X32 FILLER_0_44_193 ();
 FILLCELL_X32 FILLER_0_44_225 ();
 FILLCELL_X32 FILLER_0_44_257 ();
 FILLCELL_X32 FILLER_0_44_289 ();
 FILLCELL_X32 FILLER_0_44_321 ();
 FILLCELL_X32 FILLER_0_44_353 ();
 FILLCELL_X16 FILLER_0_44_385 ();
 FILLCELL_X8 FILLER_0_44_401 ();
 FILLCELL_X2 FILLER_0_44_409 ();
 FILLCELL_X32 FILLER_0_45_1 ();
 FILLCELL_X32 FILLER_0_45_33 ();
 FILLCELL_X32 FILLER_0_45_65 ();
 FILLCELL_X32 FILLER_0_45_97 ();
 FILLCELL_X32 FILLER_0_45_129 ();
 FILLCELL_X32 FILLER_0_45_161 ();
 FILLCELL_X32 FILLER_0_45_193 ();
 FILLCELL_X32 FILLER_0_45_225 ();
 FILLCELL_X32 FILLER_0_45_257 ();
 FILLCELL_X32 FILLER_0_45_289 ();
 FILLCELL_X32 FILLER_0_45_321 ();
 FILLCELL_X32 FILLER_0_45_353 ();
 FILLCELL_X16 FILLER_0_45_385 ();
 FILLCELL_X8 FILLER_0_45_401 ();
 FILLCELL_X2 FILLER_0_45_409 ();
 FILLCELL_X32 FILLER_0_46_1 ();
 FILLCELL_X32 FILLER_0_46_33 ();
 FILLCELL_X32 FILLER_0_46_65 ();
 FILLCELL_X32 FILLER_0_46_97 ();
 FILLCELL_X32 FILLER_0_46_129 ();
 FILLCELL_X32 FILLER_0_46_161 ();
 FILLCELL_X32 FILLER_0_46_193 ();
 FILLCELL_X32 FILLER_0_46_225 ();
 FILLCELL_X32 FILLER_0_46_257 ();
 FILLCELL_X32 FILLER_0_46_289 ();
 FILLCELL_X32 FILLER_0_46_321 ();
 FILLCELL_X32 FILLER_0_46_353 ();
 FILLCELL_X16 FILLER_0_46_385 ();
 FILLCELL_X8 FILLER_0_46_401 ();
 FILLCELL_X2 FILLER_0_46_409 ();
 FILLCELL_X32 FILLER_0_47_1 ();
 FILLCELL_X32 FILLER_0_47_33 ();
 FILLCELL_X32 FILLER_0_47_65 ();
 FILLCELL_X32 FILLER_0_47_97 ();
 FILLCELL_X32 FILLER_0_47_129 ();
 FILLCELL_X32 FILLER_0_47_161 ();
 FILLCELL_X32 FILLER_0_47_193 ();
 FILLCELL_X32 FILLER_0_47_225 ();
 FILLCELL_X32 FILLER_0_47_257 ();
 FILLCELL_X32 FILLER_0_47_289 ();
 FILLCELL_X32 FILLER_0_47_321 ();
 FILLCELL_X32 FILLER_0_47_353 ();
 FILLCELL_X16 FILLER_0_47_385 ();
 FILLCELL_X8 FILLER_0_47_401 ();
 FILLCELL_X2 FILLER_0_47_409 ();
 FILLCELL_X32 FILLER_0_48_1 ();
 FILLCELL_X32 FILLER_0_48_33 ();
 FILLCELL_X32 FILLER_0_48_65 ();
 FILLCELL_X32 FILLER_0_48_97 ();
 FILLCELL_X32 FILLER_0_48_129 ();
 FILLCELL_X32 FILLER_0_48_161 ();
 FILLCELL_X32 FILLER_0_48_193 ();
 FILLCELL_X32 FILLER_0_48_225 ();
 FILLCELL_X32 FILLER_0_48_257 ();
 FILLCELL_X32 FILLER_0_48_289 ();
 FILLCELL_X32 FILLER_0_48_321 ();
 FILLCELL_X32 FILLER_0_48_353 ();
 FILLCELL_X16 FILLER_0_48_385 ();
 FILLCELL_X8 FILLER_0_48_401 ();
 FILLCELL_X2 FILLER_0_48_409 ();
 FILLCELL_X32 FILLER_0_49_1 ();
 FILLCELL_X32 FILLER_0_49_33 ();
 FILLCELL_X32 FILLER_0_49_65 ();
 FILLCELL_X32 FILLER_0_49_97 ();
 FILLCELL_X32 FILLER_0_49_129 ();
 FILLCELL_X32 FILLER_0_49_161 ();
 FILLCELL_X32 FILLER_0_49_193 ();
 FILLCELL_X32 FILLER_0_49_225 ();
 FILLCELL_X32 FILLER_0_49_257 ();
 FILLCELL_X32 FILLER_0_49_289 ();
 FILLCELL_X32 FILLER_0_49_321 ();
 FILLCELL_X32 FILLER_0_49_353 ();
 FILLCELL_X16 FILLER_0_49_385 ();
 FILLCELL_X8 FILLER_0_49_401 ();
 FILLCELL_X2 FILLER_0_49_409 ();
 FILLCELL_X32 FILLER_0_50_1 ();
 FILLCELL_X32 FILLER_0_50_33 ();
 FILLCELL_X32 FILLER_0_50_65 ();
 FILLCELL_X32 FILLER_0_50_97 ();
 FILLCELL_X32 FILLER_0_50_129 ();
 FILLCELL_X32 FILLER_0_50_161 ();
 FILLCELL_X32 FILLER_0_50_193 ();
 FILLCELL_X32 FILLER_0_50_225 ();
 FILLCELL_X32 FILLER_0_50_257 ();
 FILLCELL_X32 FILLER_0_50_289 ();
 FILLCELL_X32 FILLER_0_50_321 ();
 FILLCELL_X32 FILLER_0_50_353 ();
 FILLCELL_X16 FILLER_0_50_385 ();
 FILLCELL_X8 FILLER_0_50_401 ();
 FILLCELL_X2 FILLER_0_50_409 ();
 FILLCELL_X32 FILLER_0_51_1 ();
 FILLCELL_X32 FILLER_0_51_33 ();
 FILLCELL_X32 FILLER_0_51_65 ();
 FILLCELL_X32 FILLER_0_51_97 ();
 FILLCELL_X32 FILLER_0_51_129 ();
 FILLCELL_X32 FILLER_0_51_161 ();
 FILLCELL_X32 FILLER_0_51_193 ();
 FILLCELL_X32 FILLER_0_51_225 ();
 FILLCELL_X32 FILLER_0_51_257 ();
 FILLCELL_X32 FILLER_0_51_289 ();
 FILLCELL_X32 FILLER_0_51_321 ();
 FILLCELL_X32 FILLER_0_51_353 ();
 FILLCELL_X16 FILLER_0_51_385 ();
 FILLCELL_X8 FILLER_0_51_401 ();
 FILLCELL_X2 FILLER_0_51_409 ();
 FILLCELL_X32 FILLER_0_52_1 ();
 FILLCELL_X32 FILLER_0_52_33 ();
 FILLCELL_X32 FILLER_0_52_65 ();
 FILLCELL_X32 FILLER_0_52_97 ();
 FILLCELL_X32 FILLER_0_52_129 ();
 FILLCELL_X32 FILLER_0_52_161 ();
 FILLCELL_X32 FILLER_0_52_193 ();
 FILLCELL_X32 FILLER_0_52_225 ();
 FILLCELL_X32 FILLER_0_52_257 ();
 FILLCELL_X32 FILLER_0_52_289 ();
 FILLCELL_X32 FILLER_0_52_321 ();
 FILLCELL_X32 FILLER_0_52_353 ();
 FILLCELL_X16 FILLER_0_52_385 ();
 FILLCELL_X8 FILLER_0_52_401 ();
 FILLCELL_X2 FILLER_0_52_409 ();
 FILLCELL_X32 FILLER_0_53_1 ();
 FILLCELL_X32 FILLER_0_53_33 ();
 FILLCELL_X32 FILLER_0_53_65 ();
 FILLCELL_X32 FILLER_0_53_97 ();
 FILLCELL_X32 FILLER_0_53_129 ();
 FILLCELL_X32 FILLER_0_53_161 ();
 FILLCELL_X32 FILLER_0_53_193 ();
 FILLCELL_X32 FILLER_0_53_225 ();
 FILLCELL_X32 FILLER_0_53_257 ();
 FILLCELL_X32 FILLER_0_53_289 ();
 FILLCELL_X32 FILLER_0_53_321 ();
 FILLCELL_X32 FILLER_0_53_353 ();
 FILLCELL_X16 FILLER_0_53_385 ();
 FILLCELL_X8 FILLER_0_53_401 ();
 FILLCELL_X2 FILLER_0_53_409 ();
 FILLCELL_X32 FILLER_0_54_1 ();
 FILLCELL_X32 FILLER_0_54_33 ();
 FILLCELL_X32 FILLER_0_54_65 ();
 FILLCELL_X32 FILLER_0_54_97 ();
 FILLCELL_X32 FILLER_0_54_129 ();
 FILLCELL_X32 FILLER_0_54_161 ();
 FILLCELL_X32 FILLER_0_54_193 ();
 FILLCELL_X32 FILLER_0_54_225 ();
 FILLCELL_X32 FILLER_0_54_257 ();
 FILLCELL_X32 FILLER_0_54_289 ();
 FILLCELL_X32 FILLER_0_54_321 ();
 FILLCELL_X32 FILLER_0_54_353 ();
 FILLCELL_X16 FILLER_0_54_385 ();
 FILLCELL_X8 FILLER_0_54_401 ();
 FILLCELL_X2 FILLER_0_54_409 ();
endmodule
