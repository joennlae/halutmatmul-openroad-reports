module fp_16_32_adder (operand_fp16_i,
    operand_fp32_i,
    result_o);
 input [15:0] operand_fp16_i;
 input [31:0] operand_fp32_i;
 output [31:0] result_o;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire net74;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire net73;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire net72;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire net71;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire net70;
 wire _0234_;
 wire net68;
 wire net67;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire net66;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire net65;
 wire net64;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire net63;
 wire net62;
 wire _0267_;
 wire net61;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire net60;
 wire _0276_;
 wire net59;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire net58;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire net57;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire net56;
 wire net55;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire net54;
 wire _0305_;
 wire net53;
 wire _0307_;
 wire _0308_;
 wire net52;
 wire net51;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire net50;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire net49;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire net48;
 wire _0336_;
 wire _0337_;
 wire net47;
 wire net46;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire net45;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire net44;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire net43;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire net42;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire net41;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire net40;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire net39;
 wire _0420_;
 wire net38;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire net37;
 wire net36;
 wire _0427_;
 wire net35;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire net34;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire net33;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire net32;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire net31;
 wire _0475_;
 wire _0476_;
 wire net30;
 wire _0478_;
 wire net29;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire net27;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire net26;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire net25;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire net24;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire net23;
 wire _0666_;
 wire net22;
 wire net21;
 wire _0669_;
 wire _0670_;
 wire net20;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire net19;
 wire _0714_;
 wire net18;
 wire _0716_;
 wire net17;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire net16;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire net15;
 wire net14;
 wire _1022_;
 wire net13;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire net12;
 wire _1049_;
 wire _1050_;
 wire net11;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire net10;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire net9;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire net8;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire net7;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire net6;
 wire net5;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire net4;
 wire _1252_;
 wire net3;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire net2;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire net1;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire net118;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire net117;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire net116;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire net114;
 wire net113;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire net112;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire net110;
 wire net109;
 wire net108;
 wire _1553_;
 wire net107;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire net105;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire net104;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire net103;
 wire net102;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire net101;
 wire _1617_;
 wire net100;
 wire net99;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire net96;
 wire net95;
 wire _1626_;
 wire _1627_;
 wire net94;
 wire net93;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire net92;
 wire _1637_;
 wire _1638_;
 wire net91;
 wire _1640_;
 wire _1641_;
 wire net90;
 wire _1643_;
 wire net89;
 wire _1645_;
 wire net88;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire net87;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire net86;
 wire net85;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire net84;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire net83;
 wire _1787_;
 wire net82;
 wire _1789_;
 wire net81;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire net80;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire net79;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire net78;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire net77;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire net76;
 wire _1897_;
 wire _1898_;
 wire net75;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire net28;
 wire _2113_;
 wire _2114_;
 wire net69;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire net115;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire net98;
 wire net97;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire net111;
 wire _2367_;
 wire _2368_;
 wire net106;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net182;
 wire net187;
 wire net192;
 wire net193;

 BUF_X1 input10 (.A(operand_fp16_i[3]),
    .Z(net10));
 NOR2_X4 _2378_ (.A1(net15),
    .A2(net16),
    .ZN(_1480_));
 NOR2_X4 _2379_ (.A1(net13),
    .A2(net14),
    .ZN(_1481_));
 NAND2_X4 _2380_ (.A1(_1481_),
    .A2(_1480_),
    .ZN(_1482_));
 BUF_X4 input9 (.A(operand_fp16_i[2]),
    .Z(net9));
 NOR2_X4 _2382_ (.A1(net11),
    .A2(net12),
    .ZN(_1484_));
 NOR2_X4 _2383_ (.A1(net10),
    .A2(net9),
    .ZN(_1485_));
 NAND2_X2 _2384_ (.A1(_1485_),
    .A2(_1484_),
    .ZN(_1486_));
 NOR2_X4 _2385_ (.A1(_1486_),
    .A2(_1482_),
    .ZN(_1487_));
 NOR2_X1 _2386_ (.A1(net5),
    .A2(net4),
    .ZN(_1488_));
 INV_X2 _2387_ (.A(net6),
    .ZN(_2195_));
 NAND2_X1 _2388_ (.A1(_1488_),
    .A2(_2195_),
    .ZN(_1489_));
 OR2_X1 _2389_ (.A1(net3),
    .A2(net2),
    .ZN(_1490_));
 NOR2_X4 _2390_ (.A1(_1489_),
    .A2(_1490_),
    .ZN(_1491_));
 BUF_X1 input8 (.A(operand_fp16_i[1]),
    .Z(net8));
 NOR2_X1 _2392_ (.A1(net8),
    .A2(net1),
    .ZN(_1493_));
 NAND3_X2 _2393_ (.A1(_1487_),
    .A2(_1491_),
    .A3(_1493_),
    .ZN(_1494_));
 NAND2_X2 _2394_ (.A1(_1494_),
    .A2(_2195_),
    .ZN(_1962_));
 INV_X1 _2395_ (.A(net1),
    .ZN(_1495_));
 OAI21_X4 _2396_ (.A(_1487_),
    .B1(net8),
    .B2(_1495_),
    .ZN(_1496_));
 INV_X1 _2397_ (.A(net16),
    .ZN(_1497_));
 INV_X1 _2398_ (.A(net14),
    .ZN(_1498_));
 OAI21_X1 _2399_ (.A(_1497_),
    .B1(_1498_),
    .B2(net15),
    .ZN(_1499_));
 INV_X1 _2400_ (.A(_1482_),
    .ZN(_1500_));
 INV_X1 _2401_ (.A(net12),
    .ZN(_1501_));
 INV_X1 _2402_ (.A(net10),
    .ZN(_1502_));
 OAI21_X1 _2403_ (.A(_1501_),
    .B1(_1502_),
    .B2(net11),
    .ZN(_1503_));
 AOI21_X2 _2404_ (.A(_1499_),
    .B1(_1500_),
    .B2(_1503_),
    .ZN(_1504_));
 NAND2_X4 _2405_ (.A1(_1504_),
    .A2(_1496_),
    .ZN(_1505_));
 BUF_X1 input7 (.A(operand_fp16_i[15]),
    .Z(net7));
 INV_X1 _2407_ (.A(_1481_),
    .ZN(_1506_));
 OAI21_X1 _2408_ (.A(_1480_),
    .B1(_1506_),
    .B2(_1484_),
    .ZN(_1507_));
 NOR2_X1 _2409_ (.A1(_1507_),
    .A2(_1487_),
    .ZN(_2227_));
 NAND2_X1 _2410_ (.A1(_1482_),
    .A2(_2218_),
    .ZN(_1508_));
 AOI21_X2 _2411_ (.A(net6),
    .B1(_1491_),
    .B2(_1508_),
    .ZN(_1954_));
 INV_X1 _2412_ (.A(_1954_),
    .ZN(_1958_));
 NAND2_X1 _2413_ (.A1(_1500_),
    .A2(_1486_),
    .ZN(_2219_));
 INV_X1 _2414_ (.A(_2219_),
    .ZN(_2237_));
 OAI21_X1 _2415_ (.A(_1487_),
    .B1(net8),
    .B2(net1),
    .ZN(_1509_));
 INV_X1 _2416_ (.A(_1509_),
    .ZN(_1510_));
 NAND2_X2 _2417_ (.A1(_2220_),
    .A2(_1510_),
    .ZN(_1511_));
 OAI21_X4 _2418_ (.A(_1511_),
    .B1(net149),
    .B2(net148),
    .ZN(_1512_));
 AOI21_X4 _2419_ (.A(net5),
    .B1(_1512_),
    .B2(_1491_),
    .ZN(_2215_));
 NAND2_X1 _2420_ (.A1(_1487_),
    .A2(_1493_),
    .ZN(_1513_));
 NAND2_X1 _2421_ (.A1(_1513_),
    .A2(_1491_),
    .ZN(_1514_));
 INV_X1 _2422_ (.A(_1514_),
    .ZN(_1515_));
 AOI21_X2 _2423_ (.A(net4),
    .B1(_1515_),
    .B2(_2221_),
    .ZN(_1946_));
 BUF_X1 input6 (.A(operand_fp16_i[14]),
    .Z(net6));
 BUF_X1 input5 (.A(operand_fp16_i[13]),
    .Z(net5));
 AOI21_X2 _2426_ (.A(net3),
    .B1(_1515_),
    .B2(_2229_),
    .ZN(_1938_));
 INV_X1 _2427_ (.A(_1505_),
    .ZN(_2226_));
 AOI21_X2 _2428_ (.A(net2),
    .B1(_2226_),
    .B2(_1491_),
    .ZN(_2270_));
 INV_X1 _2429_ (.A(_1494_),
    .ZN(_2234_));
 NAND2_X1 _2430_ (.A1(_2204_),
    .A2(_2208_),
    .ZN(_1518_));
 NAND2_X1 _2431_ (.A1(_2197_),
    .A2(_2199_),
    .ZN(_1519_));
 NOR2_X1 _2432_ (.A1(_1518_),
    .A2(_1519_),
    .ZN(_1520_));
 INV_X1 _2433_ (.A(_1520_),
    .ZN(_1521_));
 INV_X1 _2434_ (.A(_2216_),
    .ZN(_1522_));
 INV_X1 _2435_ (.A(_2214_),
    .ZN(_1523_));
 INV_X1 _2436_ (.A(_2224_),
    .ZN(_1524_));
 OAI21_X1 _2437_ (.A(_1522_),
    .B1(_1523_),
    .B2(_1524_),
    .ZN(_1525_));
 INV_X2 _2438_ (.A(_1525_),
    .ZN(_1526_));
 NAND2_X1 _2439_ (.A1(_2223_),
    .A2(_2214_),
    .ZN(_1527_));
 OR2_X4 _2440_ (.A1(_1944_),
    .A2(_1527_),
    .ZN(_1528_));
 AOI21_X4 _2441_ (.A(_1521_),
    .B1(_1526_),
    .B2(_1528_),
    .ZN(_1529_));
 INV_X1 _2442_ (.A(_2205_),
    .ZN(_1530_));
 INV_X1 _2443_ (.A(_2204_),
    .ZN(_1531_));
 INV_X1 _2444_ (.A(_2209_),
    .ZN(_1532_));
 OAI21_X1 _2445_ (.A(_1530_),
    .B1(_1531_),
    .B2(_1532_),
    .ZN(_1533_));
 INV_X1 _2446_ (.A(_1519_),
    .ZN(_1534_));
 NAND2_X1 _2447_ (.A1(_1533_),
    .A2(_1534_),
    .ZN(_1535_));
 INV_X1 _2448_ (.A(_2196_),
    .ZN(_1536_));
 INV_X1 _2449_ (.A(_2197_),
    .ZN(_1537_));
 INV_X1 _2450_ (.A(_2200_),
    .ZN(_1538_));
 OAI21_X1 _2451_ (.A(_1536_),
    .B1(_1537_),
    .B2(_1538_),
    .ZN(_1539_));
 INV_X1 _2452_ (.A(_1539_),
    .ZN(_1540_));
 NAND2_X1 _2453_ (.A1(_1535_),
    .A2(_1540_),
    .ZN(_1541_));
 NOR2_X4 _2454_ (.A1(_1541_),
    .A2(_1529_),
    .ZN(_1542_));
 BUF_X1 input4 (.A(operand_fp16_i[12]),
    .Z(net4));
 NAND2_X1 _2456_ (.A1(_1542_),
    .A2(_1940_),
    .ZN(_1544_));
 INV_X1 _2457_ (.A(_1945_),
    .ZN(_1545_));
 OAI21_X4 _2458_ (.A(_1544_),
    .B1(_1545_),
    .B2(net112),
    .ZN(_1546_));
 BUF_X1 input3 (.A(operand_fp16_i[11]),
    .Z(net3));
 INV_X1 _2460_ (.A(_1541_),
    .ZN(_1547_));
 NAND2_X2 _2461_ (.A1(_1526_),
    .A2(_1528_),
    .ZN(_1959_));
 NAND2_X1 _2462_ (.A1(_1959_),
    .A2(_1520_),
    .ZN(_1548_));
 NAND2_X4 _2463_ (.A1(_1548_),
    .A2(_1547_),
    .ZN(_1549_));
 BUF_X1 input2 (.A(operand_fp16_i[10]),
    .Z(net2));
 BUF_X1 input1 (.A(operand_fp16_i[0]),
    .Z(net1));
 TAPCELL_X1 PHY_109 ();
 MUX2_X2 _2467_ (.A(_1948_),
    .B(_1952_),
    .S(_1549_),
    .Z(_1553_));
 TAPCELL_X1 PHY_108 ();
 TAPCELL_X1 PHY_107 ();
 NAND2_X1 _2470_ (.A1(net90),
    .A2(_1957_),
    .ZN(_1555_));
 NAND2_X1 _2471_ (.A1(net124),
    .A2(_1961_),
    .ZN(_1556_));
 AND2_X2 _2472_ (.A1(_1555_),
    .A2(_1556_),
    .ZN(_2374_));
 INV_X1 _2473_ (.A(_2203_),
    .ZN(_1557_));
 INV_X1 _2474_ (.A(_2207_),
    .ZN(_1558_));
 OAI21_X1 _2475_ (.A(_1557_),
    .B1(_1531_),
    .B2(_1558_),
    .ZN(_1559_));
 INV_X1 _2476_ (.A(_2213_),
    .ZN(_1560_));
 INV_X1 _2477_ (.A(_2222_),
    .ZN(_1561_));
 OAI221_X2 _2478_ (.A(_1560_),
    .B1(_1523_),
    .B2(_1561_),
    .C1(_1939_),
    .C2(_1527_),
    .ZN(_1955_));
 INV_X1 _2479_ (.A(_1518_),
    .ZN(_1562_));
 AOI21_X1 _2480_ (.A(_1559_),
    .B1(_1955_),
    .B2(_1562_),
    .ZN(_1963_));
 AOI21_X1 _2481_ (.A(_1533_),
    .B1(_1959_),
    .B2(_1562_),
    .ZN(_1968_));
 MUX2_X2 _2482_ (.A(_1965_),
    .B(_1970_),
    .S(net124),
    .Z(_2357_));
 MUX2_X1 _2483_ (.A(_1956_),
    .B(_1960_),
    .S(_1549_),
    .Z(_1563_));
 XNOR2_X2 _2484_ (.A(_1531_),
    .B(_1563_),
    .ZN(_1564_));
 NOR2_X4 _2485_ (.A1(_1564_),
    .A2(_2374_),
    .ZN(_1565_));
 XNOR2_X1 _2486_ (.A(_1537_),
    .B(_1969_),
    .ZN(_1566_));
 NAND2_X1 _2487_ (.A1(net124),
    .A2(_1566_),
    .ZN(_1567_));
 XNOR2_X1 _2488_ (.A(_2197_),
    .B(_1964_),
    .ZN(_1568_));
 OAI21_X2 _2489_ (.A(_1567_),
    .B1(net124),
    .B2(_1568_),
    .ZN(_1569_));
 NAND2_X4 _2490_ (.A1(_2357_),
    .A2(_1569_),
    .ZN(_1570_));
 INV_X4 _2491_ (.A(_1570_),
    .ZN(_1571_));
 TAPCELL_X1 PHY_106 ();
 OR2_X1 _2493_ (.A1(_1549_),
    .A2(_1947_),
    .ZN(_1573_));
 OAI21_X1 _2494_ (.A(_1573_),
    .B1(_1951_),
    .B2(_1542_),
    .ZN(_1574_));
 XNOR2_X2 _2495_ (.A(net108),
    .B(_1574_),
    .ZN(_1575_));
 INV_X8 _2496_ (.A(_1553_),
    .ZN(_1576_));
 INV_X1 _2497_ (.A(_2367_),
    .ZN(_1577_));
 NOR3_X1 _2498_ (.A1(_1576_),
    .A2(_2235_),
    .A3(_1577_),
    .ZN(_1578_));
 NAND4_X1 _2499_ (.A1(_1565_),
    .A2(_1571_),
    .A3(_1575_),
    .A4(_1578_),
    .ZN(_1579_));
 NOR2_X1 _2500_ (.A1(net116),
    .A2(_1495_),
    .ZN(_1580_));
 INV_X1 _2501_ (.A(_1580_),
    .ZN(_1581_));
 TAPCELL_X1 PHY_105 ();
 NOR3_X1 _2503_ (.A1(_1581_),
    .A2(net125),
    .A3(_2239_),
    .ZN(_1583_));
 XNOR2_X2 _2504_ (.A(_1509_),
    .B(_2238_),
    .ZN(_1584_));
 NOR2_X2 _2505_ (.A1(_1584_),
    .A2(_1514_),
    .ZN(_1585_));
 INV_X2 _2506_ (.A(_1491_),
    .ZN(_1586_));
 AOI22_X2 _2507_ (.A1(_1583_),
    .A2(_1585_),
    .B1(net1),
    .B2(_1586_),
    .ZN(_1587_));
 OAI21_X1 _2508_ (.A(_2266_),
    .B1(_1587_),
    .B2(net21),
    .ZN(_1588_));
 INV_X1 _2509_ (.A(_2265_),
    .ZN(_1589_));
 NAND2_X1 _2510_ (.A1(_1588_),
    .A2(_1589_),
    .ZN(_1590_));
 NAND3_X1 _2511_ (.A1(_1590_),
    .A2(_2260_),
    .A3(_2263_),
    .ZN(_1591_));
 INV_X1 _2512_ (.A(_2259_),
    .ZN(_1592_));
 NAND2_X1 _2513_ (.A1(_2260_),
    .A2(_2262_),
    .ZN(_1593_));
 NAND3_X1 _2514_ (.A1(_1591_),
    .A2(_1592_),
    .A3(_1593_),
    .ZN(_1594_));
 NAND2_X1 _2515_ (.A1(_2248_),
    .A2(_2251_),
    .ZN(_1595_));
 INV_X1 _2516_ (.A(_1595_),
    .ZN(_1596_));
 NAND4_X1 _2517_ (.A1(_1594_),
    .A2(_2254_),
    .A3(_2257_),
    .A4(_1596_),
    .ZN(_1597_));
 NAND2_X1 _2518_ (.A1(_2256_),
    .A2(_2254_),
    .ZN(_1598_));
 INV_X1 _2519_ (.A(_1598_),
    .ZN(_1599_));
 OAI21_X1 _2520_ (.A(_1596_),
    .B1(_1599_),
    .B2(_2253_),
    .ZN(_1600_));
 INV_X1 _2521_ (.A(_2247_),
    .ZN(_1601_));
 NAND2_X1 _2522_ (.A1(_2248_),
    .A2(_2250_),
    .ZN(_1602_));
 NAND3_X1 _2523_ (.A1(_1600_),
    .A2(_1601_),
    .A3(_1602_),
    .ZN(_1603_));
 INV_X1 _2524_ (.A(_1603_),
    .ZN(_1604_));
 NAND2_X1 _2525_ (.A1(_1597_),
    .A2(_1604_),
    .ZN(_1605_));
 NAND3_X1 _2526_ (.A1(_1605_),
    .A2(_2242_),
    .A3(_2245_),
    .ZN(_1606_));
 INV_X1 _2527_ (.A(_2241_),
    .ZN(_1607_));
 NAND2_X1 _2528_ (.A1(_2242_),
    .A2(_2244_),
    .ZN(_1608_));
 NAND3_X1 _2529_ (.A1(_1606_),
    .A2(_1607_),
    .A3(_1608_),
    .ZN(_1609_));
 AOI21_X2 _2530_ (.A(_1579_),
    .B1(_1609_),
    .B2(_2236_),
    .ZN(_1610_));
 TAPCELL_X1 PHY_104 ();
 TAPCELL_X1 PHY_103 ();
 NOR2_X1 _2533_ (.A1(_1610_),
    .A2(net90),
    .ZN(_1613_));
 NAND2_X1 _2534_ (.A1(_1613_),
    .A2(net41),
    .ZN(_1614_));
 INV_X1 _2535_ (.A(net7),
    .ZN(_1615_));
 OAI21_X1 _2536_ (.A(_1614_),
    .B1(_1615_),
    .B2(_1613_),
    .ZN(net73));
 TAPCELL_X1 PHY_102 ();
 INV_X8 _2538_ (.A(net92),
    .ZN(_1617_));
 TAPCELL_X1 PHY_101 ();
 TAPCELL_X1 PHY_100 ();
 TAPCELL_X1 PHY_99 ();
 INV_X8 _2542_ (.A(_1546_),
    .ZN(_1620_));
 TAPCELL_X1 PHY_98 ();
 INV_X1 _2544_ (.A(net41),
    .ZN(_1621_));
 NAND2_X2 _2545_ (.A1(_1621_),
    .A2(net7),
    .ZN(_1622_));
 NAND2_X2 _2546_ (.A1(_1615_),
    .A2(net41),
    .ZN(_1623_));
 NAND2_X4 _2547_ (.A1(_1622_),
    .A2(_1623_),
    .ZN(_2040_));
 TAPCELL_X1 PHY_97 ();
 TAPCELL_X1 PHY_96 ();
 NAND2_X1 _2550_ (.A1(_1610_),
    .A2(net101),
    .ZN(_1626_));
 NAND2_X4 _2551_ (.A1(_1626_),
    .A2(_2040_),
    .ZN(_1627_));
 TAPCELL_X1 PHY_95 ();
 TAPCELL_X1 PHY_94 ();
 NAND2_X1 _2554_ (.A1(net101),
    .A2(_2234_),
    .ZN(_1630_));
 NOR4_X1 _2555_ (.A1(net37),
    .A2(net36),
    .A3(net40),
    .A4(net38),
    .ZN(_1631_));
 NOR4_X1 _2556_ (.A1(net33),
    .A2(net32),
    .A3(net35),
    .A4(net34),
    .ZN(_1632_));
 NAND2_X1 _2557_ (.A1(_1631_),
    .A2(_1632_),
    .ZN(_2233_));
 OAI21_X2 _2558_ (.A(_1630_),
    .B1(_2233_),
    .B2(net101),
    .ZN(_1633_));
 NOR3_X1 _2559_ (.A1(_1570_),
    .A2(_1617_),
    .A3(_1633_),
    .ZN(_1634_));
 INV_X1 _2560_ (.A(_1634_),
    .ZN(_1635_));
 TAPCELL_X1 PHY_93 ();
 NOR2_X1 _2562_ (.A1(_1635_),
    .A2(net129),
    .ZN(_1637_));
 INV_X1 _2563_ (.A(_1637_),
    .ZN(_1638_));
 TAPCELL_X1 PHY_92 ();
 NOR2_X1 _2565_ (.A1(_1638_),
    .A2(_1576_),
    .ZN(_1640_));
 INV_X1 _2566_ (.A(_1640_),
    .ZN(_1641_));
 TAPCELL_X1 PHY_91 ();
 INV_X4 _2568_ (.A(net97),
    .ZN(_1643_));
 TAPCELL_X1 PHY_90 ();
 NOR2_X1 _2570_ (.A1(_1641_),
    .A2(_1643_),
    .ZN(_1645_));
 TAPCELL_X1 PHY_89 ();
 NAND2_X1 _2572_ (.A1(_1645_),
    .A2(_1565_),
    .ZN(_1647_));
 XNOR2_X1 _2573_ (.A(_1627_),
    .B(_1647_),
    .ZN(_1973_));
 NAND3_X4 _2574_ (.A1(_1610_),
    .A2(net101),
    .A3(_2040_),
    .ZN(_1648_));
 INV_X2 _2575_ (.A(_1648_),
    .ZN(_2033_));
 NAND2_X1 _2576_ (.A1(_2233_),
    .A2(net101),
    .ZN(_1649_));
 OAI21_X1 _2577_ (.A(_1649_),
    .B1(_2234_),
    .B2(net101),
    .ZN(_1650_));
 XNOR2_X1 _2578_ (.A(_2033_),
    .B(_1650_),
    .ZN(_1972_));
 NAND2_X1 _2579_ (.A1(_1586_),
    .A2(net16),
    .ZN(_1651_));
 INV_X1 _2580_ (.A(net11),
    .ZN(_1652_));
 NAND2_X1 _2581_ (.A1(_1505_),
    .A2(_1652_),
    .ZN(_1653_));
 OAI21_X1 _2582_ (.A(_1653_),
    .B1(net12),
    .B2(net116),
    .ZN(_1654_));
 INV_X2 _2583_ (.A(net96),
    .ZN(_1655_));
 NAND2_X1 _2584_ (.A1(_1654_),
    .A2(_1655_),
    .ZN(_1656_));
 INV_X1 _2585_ (.A(net9),
    .ZN(_1657_));
 NAND2_X1 _2586_ (.A1(_1505_),
    .A2(_1657_),
    .ZN(_1658_));
 OAI21_X1 _2587_ (.A(_1658_),
    .B1(net10),
    .B2(net116),
    .ZN(_1659_));
 INV_X1 _2588_ (.A(_1659_),
    .ZN(_1660_));
 OAI21_X1 _2589_ (.A(_1656_),
    .B1(_1655_),
    .B2(_1660_),
    .ZN(_1661_));
 NAND2_X1 _2590_ (.A1(_1661_),
    .A2(_2239_),
    .ZN(_1662_));
 INV_X2 _2591_ (.A(_2239_),
    .ZN(_1663_));
 NAND2_X1 _2592_ (.A1(net116),
    .A2(net13),
    .ZN(_1664_));
 OAI21_X1 _2593_ (.A(_1664_),
    .B1(_1498_),
    .B2(net121),
    .ZN(_1665_));
 NOR2_X1 _2594_ (.A1(_1665_),
    .A2(_1655_),
    .ZN(_1666_));
 AOI21_X1 _2595_ (.A(net96),
    .B1(net116),
    .B2(net15),
    .ZN(_1667_));
 OAI21_X1 _2596_ (.A(_1663_),
    .B1(_1666_),
    .B2(_1667_),
    .ZN(_1668_));
 AOI21_X1 _2597_ (.A(_1584_),
    .B1(_1662_),
    .B2(_1668_),
    .ZN(_1669_));
 NAND2_X1 _2598_ (.A1(_1505_),
    .A2(_1495_),
    .ZN(_1670_));
 OAI21_X1 _2599_ (.A(_1670_),
    .B1(net8),
    .B2(net121),
    .ZN(_1671_));
 NOR2_X1 _2600_ (.A1(_1671_),
    .A2(net96),
    .ZN(_1672_));
 NAND2_X1 _2601_ (.A1(_1672_),
    .A2(_1663_),
    .ZN(_1673_));
 INV_X1 _2602_ (.A(_1673_),
    .ZN(_1674_));
 INV_X1 _2603_ (.A(_1584_),
    .ZN(_1675_));
 OAI21_X1 _2604_ (.A(_1515_),
    .B1(_1674_),
    .B2(_1675_),
    .ZN(_1676_));
 OAI21_X1 _2605_ (.A(_1651_),
    .B1(_1669_),
    .B2(_1676_),
    .ZN(_1677_));
 INV_X1 _2606_ (.A(_1677_),
    .ZN(_2240_));
 NAND2_X1 _2607_ (.A1(net121),
    .A2(_1502_),
    .ZN(_1678_));
 OAI21_X1 _2608_ (.A(_1678_),
    .B1(net11),
    .B2(net116),
    .ZN(_1679_));
 NAND2_X1 _2609_ (.A1(_1679_),
    .A2(_1655_),
    .ZN(_1680_));
 INV_X1 _2610_ (.A(net8),
    .ZN(_1681_));
 NAND2_X1 _2611_ (.A1(net121),
    .A2(_1681_),
    .ZN(_1682_));
 OAI21_X1 _2612_ (.A(_1682_),
    .B1(net9),
    .B2(net116),
    .ZN(_1683_));
 INV_X1 _2613_ (.A(_1683_),
    .ZN(_1684_));
 OAI21_X1 _2614_ (.A(_1680_),
    .B1(_1655_),
    .B2(_1684_),
    .ZN(_1685_));
 AND2_X1 _2615_ (.A1(_1685_),
    .A2(_2239_),
    .ZN(_1686_));
 NAND2_X1 _2616_ (.A1(net121),
    .A2(_1501_),
    .ZN(_1687_));
 OAI21_X1 _2617_ (.A(_1687_),
    .B1(net13),
    .B2(net116),
    .ZN(_1688_));
 NAND2_X1 _2618_ (.A1(_1688_),
    .A2(net125),
    .ZN(_1689_));
 NOR2_X1 _2619_ (.A1(_2226_),
    .A2(net14),
    .ZN(_1690_));
 NOR2_X1 _2620_ (.A1(net116),
    .A2(net15),
    .ZN(_1691_));
 OAI21_X1 _2621_ (.A(_1655_),
    .B1(_1690_),
    .B2(_1691_),
    .ZN(_1692_));
 AOI21_X1 _2622_ (.A(_2239_),
    .B1(_1689_),
    .B2(_1692_),
    .ZN(_1693_));
 OAI21_X1 _2623_ (.A(_1675_),
    .B1(_1686_),
    .B2(_1693_),
    .ZN(_1694_));
 INV_X1 _2624_ (.A(_1583_),
    .ZN(_1695_));
 AOI21_X1 _2625_ (.A(_1514_),
    .B1(_1695_),
    .B2(_1584_),
    .ZN(_1696_));
 NAND2_X1 _2626_ (.A1(_1694_),
    .A2(_1696_),
    .ZN(_1697_));
 NAND2_X1 _2627_ (.A1(_1586_),
    .A2(net15),
    .ZN(_1698_));
 NAND2_X1 _2628_ (.A1(_1697_),
    .A2(_1698_),
    .ZN(_1699_));
 INV_X1 _2629_ (.A(_1699_),
    .ZN(_2243_));
 INV_X1 _2630_ (.A(_1585_),
    .ZN(_1700_));
 NAND2_X1 _2631_ (.A1(_1654_),
    .A2(net96),
    .ZN(_1701_));
 OAI21_X1 _2632_ (.A(_1701_),
    .B1(net96),
    .B2(_1665_),
    .ZN(_1702_));
 AOI21_X1 _2633_ (.A(_1700_),
    .B1(_1702_),
    .B2(_1663_),
    .ZN(_1703_));
 NAND2_X1 _2634_ (.A1(_1660_),
    .A2(_1655_),
    .ZN(_1704_));
 OAI21_X1 _2635_ (.A(_1704_),
    .B1(_1655_),
    .B2(_1671_),
    .ZN(_1705_));
 OAI21_X1 _2636_ (.A(_1703_),
    .B1(_1663_),
    .B2(_1705_),
    .ZN(_1706_));
 NAND2_X1 _2637_ (.A1(_1586_),
    .A2(net14),
    .ZN(_1707_));
 NAND2_X1 _2638_ (.A1(_1706_),
    .A2(_1707_),
    .ZN(_1708_));
 INV_X1 _2639_ (.A(_1708_),
    .ZN(_2246_));
 NAND2_X1 _2640_ (.A1(_1679_),
    .A2(net96),
    .ZN(_1709_));
 INV_X1 _2641_ (.A(_1688_),
    .ZN(_1710_));
 OAI21_X1 _2642_ (.A(_1709_),
    .B1(net96),
    .B2(_1710_),
    .ZN(_1711_));
 AOI21_X1 _2643_ (.A(_1700_),
    .B1(_1711_),
    .B2(_1663_),
    .ZN(_1712_));
 NAND2_X1 _2644_ (.A1(_1580_),
    .A2(net96),
    .ZN(_1713_));
 OAI21_X2 _2645_ (.A(_1713_),
    .B1(_1683_),
    .B2(net96),
    .ZN(_1714_));
 OAI21_X1 _2646_ (.A(_1712_),
    .B1(_1663_),
    .B2(_1714_),
    .ZN(_1715_));
 NAND2_X1 _2647_ (.A1(_1586_),
    .A2(net13),
    .ZN(_1716_));
 NAND2_X1 _2648_ (.A1(_1715_),
    .A2(_1716_),
    .ZN(_1717_));
 INV_X1 _2649_ (.A(_1717_),
    .ZN(_2249_));
 NAND2_X1 _2650_ (.A1(_1661_),
    .A2(_1663_),
    .ZN(_1718_));
 OAI21_X1 _2651_ (.A(_2239_),
    .B1(_1671_),
    .B2(net126),
    .ZN(_1719_));
 NAND3_X1 _2652_ (.A1(_1718_),
    .A2(_1585_),
    .A3(_1719_),
    .ZN(_1720_));
 OAI21_X1 _2653_ (.A(_1720_),
    .B1(_1501_),
    .B2(_1491_),
    .ZN(_1721_));
 INV_X1 _2654_ (.A(_1721_),
    .ZN(_2252_));
 NAND2_X1 _2655_ (.A1(_1685_),
    .A2(_1663_),
    .ZN(_1722_));
 OAI21_X1 _2656_ (.A(_2239_),
    .B1(_1581_),
    .B2(net126),
    .ZN(_1723_));
 NAND3_X1 _2657_ (.A1(_1722_),
    .A2(_1585_),
    .A3(_1723_),
    .ZN(_1724_));
 NAND2_X1 _2658_ (.A1(_1586_),
    .A2(net11),
    .ZN(_1725_));
 NAND2_X1 _2659_ (.A1(_1724_),
    .A2(_1725_),
    .ZN(_1726_));
 INV_X1 _2660_ (.A(_1726_),
    .ZN(_2255_));
 NAND2_X1 _2661_ (.A1(_1585_),
    .A2(_1663_),
    .ZN(_1727_));
 INV_X1 _2662_ (.A(_1727_),
    .ZN(_1728_));
 NAND2_X1 _2663_ (.A1(_1705_),
    .A2(_1728_),
    .ZN(_1729_));
 NAND2_X1 _2664_ (.A1(_1586_),
    .A2(net10),
    .ZN(_1730_));
 NAND2_X1 _2665_ (.A1(_1729_),
    .A2(_1730_),
    .ZN(_1731_));
 INV_X1 _2666_ (.A(_1731_),
    .ZN(_2258_));
 AOI22_X4 _2667_ (.A1(_1714_),
    .A2(_1728_),
    .B1(net9),
    .B2(_1586_),
    .ZN(_2261_));
 OAI22_X1 _2668_ (.A1(_1673_),
    .A2(_1700_),
    .B1(_1681_),
    .B2(_1491_),
    .ZN(_1732_));
 INV_X1 _2669_ (.A(_1732_),
    .ZN(_2264_));
 INV_X4 _2670_ (.A(_1627_),
    .ZN(_1733_));
 NAND2_X1 _2671_ (.A1(_2264_),
    .A2(net109),
    .ZN(_1734_));
 TAPCELL_X1 PHY_88 ();
 OR2_X1 _2673_ (.A1(net109),
    .A2(net22),
    .ZN(_1736_));
 NAND3_X1 _2674_ (.A1(_1734_),
    .A2(_1571_),
    .A3(_1736_),
    .ZN(_1737_));
 NAND2_X1 _2675_ (.A1(_1737_),
    .A2(_1617_),
    .ZN(_1738_));
 OR2_X1 _2676_ (.A1(net109),
    .A2(net21),
    .ZN(_1739_));
 INV_X1 _2677_ (.A(_1587_),
    .ZN(_1740_));
 OAI21_X1 _2678_ (.A(_1739_),
    .B1(_1740_),
    .B2(net90),
    .ZN(_1741_));
 INV_X1 _2679_ (.A(_1741_),
    .ZN(_1742_));
 NAND2_X1 _2680_ (.A1(_1742_),
    .A2(_1571_),
    .ZN(_1743_));
 INV_X1 _2681_ (.A(_1743_),
    .ZN(_1744_));
 OAI21_X1 _2682_ (.A(_1738_),
    .B1(_1617_),
    .B2(_1744_),
    .ZN(_1745_));
 NAND2_X1 _2683_ (.A1(_2261_),
    .A2(net109),
    .ZN(_1746_));
 OR2_X1 _2684_ (.A1(net109),
    .A2(net23),
    .ZN(_1747_));
 NAND2_X1 _2685_ (.A1(_1746_),
    .A2(_1747_),
    .ZN(_1748_));
 INV_X1 _2686_ (.A(_1748_),
    .ZN(_1749_));
 NAND2_X1 _2687_ (.A1(_1749_),
    .A2(_1571_),
    .ZN(_1750_));
 TAPCELL_X1 PHY_87 ();
 TAPCELL_X1 PHY_86 ();
 NAND2_X1 _2690_ (.A1(_1750_),
    .A2(net94),
    .ZN(_1753_));
 NOR2_X1 _2691_ (.A1(net109),
    .A2(net24),
    .ZN(_1754_));
 AOI21_X2 _2692_ (.A(_1754_),
    .B1(_2258_),
    .B2(net101),
    .ZN(_1755_));
 NAND2_X1 _2693_ (.A1(_1755_),
    .A2(_1571_),
    .ZN(_1756_));
 INV_X1 _2694_ (.A(_1756_),
    .ZN(_1757_));
 OAI21_X1 _2695_ (.A(_1753_),
    .B1(_1757_),
    .B2(net94),
    .ZN(_1758_));
 MUX2_X1 _2696_ (.A(_1745_),
    .B(_1758_),
    .S(_1620_),
    .Z(_1759_));
 INV_X1 _2697_ (.A(_1759_),
    .ZN(_1760_));
 NOR2_X1 _2698_ (.A1(_1760_),
    .A2(_1576_),
    .ZN(_1761_));
 OR2_X1 _2699_ (.A1(net101),
    .A2(net25),
    .ZN(_1762_));
 OAI21_X1 _2700_ (.A(_1762_),
    .B1(_1726_),
    .B2(net90),
    .ZN(_1763_));
 INV_X1 _2701_ (.A(_1763_),
    .ZN(_1764_));
 NAND2_X1 _2702_ (.A1(_1764_),
    .A2(_1571_),
    .ZN(_1765_));
 NAND2_X1 _2703_ (.A1(_1765_),
    .A2(net94),
    .ZN(_1766_));
 OR2_X1 _2704_ (.A1(net101),
    .A2(net26),
    .ZN(_1767_));
 OAI21_X1 _2705_ (.A(_1767_),
    .B1(_1721_),
    .B2(net90),
    .ZN(_1768_));
 INV_X1 _2706_ (.A(_1768_),
    .ZN(_1769_));
 NAND2_X1 _2707_ (.A1(_1769_),
    .A2(_1571_),
    .ZN(_1770_));
 INV_X1 _2708_ (.A(_1770_),
    .ZN(_1771_));
 TAPCELL_X1 PHY_85 ();
 OAI21_X1 _2710_ (.A(_1766_),
    .B1(_1771_),
    .B2(net94),
    .ZN(_1773_));
 NAND2_X1 _2711_ (.A1(_1773_),
    .A2(net110),
    .ZN(_1774_));
 NAND2_X1 _2712_ (.A1(_2249_),
    .A2(net109),
    .ZN(_1775_));
 OR2_X1 _2713_ (.A1(net101),
    .A2(net27),
    .ZN(_1776_));
 NAND2_X1 _2714_ (.A1(_1775_),
    .A2(_1776_),
    .ZN(_1777_));
 INV_X1 _2715_ (.A(_1777_),
    .ZN(_1778_));
 NAND3_X1 _2716_ (.A1(_1778_),
    .A2(net95),
    .A3(_1571_),
    .ZN(_1779_));
 NAND2_X1 _2717_ (.A1(_2246_),
    .A2(net101),
    .ZN(_1780_));
 OAI21_X1 _2718_ (.A(_1780_),
    .B1(net29),
    .B2(net101),
    .ZN(_1781_));
 INV_X1 _2719_ (.A(_1781_),
    .ZN(_1782_));
 NAND2_X1 _2720_ (.A1(_1782_),
    .A2(_1571_),
    .ZN(_1783_));
 OAI21_X1 _2721_ (.A(_1779_),
    .B1(_1783_),
    .B2(net95),
    .ZN(_1784_));
 OAI21_X1 _2722_ (.A(_1774_),
    .B1(_1784_),
    .B2(net110),
    .ZN(_1785_));
 TAPCELL_X1 PHY_84 ();
 AOI21_X1 _2724_ (.A(_1761_),
    .B1(_1785_),
    .B2(_1576_),
    .ZN(_1787_));
 TAPCELL_X1 PHY_83 ();
 NAND2_X1 _2726_ (.A1(_1787_),
    .A2(net89),
    .ZN(_1789_));
 TAPCELL_X1 PHY_82 ();
 NAND2_X1 _2728_ (.A1(_2240_),
    .A2(net101),
    .ZN(_1791_));
 OR2_X1 _2729_ (.A1(net101),
    .A2(net31),
    .ZN(_1792_));
 NAND3_X1 _2730_ (.A1(_1791_),
    .A2(_1571_),
    .A3(_1792_),
    .ZN(_1793_));
 TAPCELL_X1 PHY_81 ();
 NAND2_X1 _2732_ (.A1(_1793_),
    .A2(_1617_),
    .ZN(_1795_));
 NAND3_X1 _2733_ (.A1(_1697_),
    .A2(net101),
    .A3(_1698_),
    .ZN(_1796_));
 OR2_X1 _2734_ (.A1(net101),
    .A2(net30),
    .ZN(_1797_));
 NAND2_X1 _2735_ (.A1(_1796_),
    .A2(_1797_),
    .ZN(_1798_));
 INV_X1 _2736_ (.A(_1798_),
    .ZN(_1799_));
 NAND2_X1 _2737_ (.A1(_1799_),
    .A2(_1571_),
    .ZN(_1800_));
 INV_X1 _2738_ (.A(_1800_),
    .ZN(_1801_));
 OAI21_X1 _2739_ (.A(_1795_),
    .B1(_1801_),
    .B2(_1617_),
    .ZN(_1802_));
 NAND2_X1 _2740_ (.A1(_1802_),
    .A2(net110),
    .ZN(_1803_));
 OAI21_X1 _2741_ (.A(_1803_),
    .B1(net110),
    .B2(_1634_),
    .ZN(_1804_));
 NOR2_X1 _2742_ (.A1(_1804_),
    .A2(_1576_),
    .ZN(_1805_));
 INV_X1 _2743_ (.A(_1805_),
    .ZN(_1806_));
 OAI21_X1 _2744_ (.A(_1789_),
    .B1(net97),
    .B2(_1806_),
    .ZN(_1807_));
 NAND3_X1 _2745_ (.A1(_1733_),
    .A2(_1565_),
    .A3(_1807_),
    .ZN(_1808_));
 NAND2_X1 _2746_ (.A1(_1807_),
    .A2(_1565_),
    .ZN(_1809_));
 NAND2_X1 _2747_ (.A1(_1809_),
    .A2(_1627_),
    .ZN(_1810_));
 NAND2_X1 _2748_ (.A1(_1808_),
    .A2(_1810_),
    .ZN(_1998_));
 NOR2_X1 _2749_ (.A1(net90),
    .A2(net21),
    .ZN(_1811_));
 TAPCELL_X1 PHY_80 ();
 AOI21_X1 _2751_ (.A(_1811_),
    .B1(_1587_),
    .B2(net90),
    .ZN(_1813_));
 XNOR2_X1 _2752_ (.A(_2033_),
    .B(_1813_),
    .ZN(_1997_));
 INV_X2 _2753_ (.A(_1565_),
    .ZN(_1814_));
 INV_X1 _2754_ (.A(net18),
    .ZN(_1815_));
 NOR2_X1 _2755_ (.A1(net123),
    .A2(_1815_),
    .ZN(_1816_));
 INV_X1 _2756_ (.A(_1816_),
    .ZN(_1817_));
 OAI21_X1 _2757_ (.A(_1617_),
    .B1(_1570_),
    .B2(_1817_),
    .ZN(_1818_));
 INV_X1 _2758_ (.A(net48),
    .ZN(_1819_));
 NOR2_X1 _2759_ (.A1(net109),
    .A2(_1819_),
    .ZN(_1820_));
 AND2_X1 _2760_ (.A1(_1571_),
    .A2(_1820_),
    .ZN(_1821_));
 OAI21_X1 _2761_ (.A(_1818_),
    .B1(_1821_),
    .B2(_1617_),
    .ZN(_1822_));
 INV_X1 _2762_ (.A(net20),
    .ZN(_1823_));
 NOR2_X1 _2763_ (.A1(net123),
    .A2(_1823_),
    .ZN(_1824_));
 NAND2_X1 _2764_ (.A1(_1571_),
    .A2(_1824_),
    .ZN(_1825_));
 INV_X1 _2765_ (.A(net19),
    .ZN(_1826_));
 NOR2_X1 _2766_ (.A1(net109),
    .A2(_1826_),
    .ZN(_1827_));
 NAND2_X1 _2767_ (.A1(_1571_),
    .A2(_1827_),
    .ZN(_1828_));
 MUX2_X1 _2768_ (.A(_1825_),
    .B(_1828_),
    .S(net93),
    .Z(_1829_));
 MUX2_X1 _2769_ (.A(_1822_),
    .B(_1829_),
    .S(net145),
    .Z(_1830_));
 NOR2_X1 _2770_ (.A1(_1830_),
    .A2(_1576_),
    .ZN(_1831_));
 AOI21_X1 _2771_ (.A(_1831_),
    .B1(_1760_),
    .B2(_1576_),
    .ZN(_1832_));
 AOI21_X1 _2772_ (.A(_1814_),
    .B1(_1832_),
    .B2(net89),
    .ZN(_1833_));
 OR2_X1 _2773_ (.A1(_1804_),
    .A2(net105),
    .ZN(_1834_));
 OR2_X1 _2774_ (.A1(_1785_),
    .A2(_1576_),
    .ZN(_1835_));
 NAND2_X1 _2775_ (.A1(_1834_),
    .A2(_1835_),
    .ZN(_1836_));
 OAI21_X1 _2776_ (.A(_1833_),
    .B1(_1836_),
    .B2(net89),
    .ZN(_1837_));
 OR2_X1 _2777_ (.A1(_1627_),
    .A2(_1837_),
    .ZN(_1838_));
 NAND2_X1 _2778_ (.A1(_1627_),
    .A2(_1837_),
    .ZN(_1839_));
 NAND2_X1 _2779_ (.A1(_1838_),
    .A2(_1839_),
    .ZN(_2008_));
 TAPCELL_X1 PHY_79 ();
 NAND2_X1 _2781_ (.A1(net101),
    .A2(net48),
    .ZN(_1841_));
 XNOR2_X2 _2782_ (.A(_1648_),
    .B(_1841_),
    .ZN(_2007_));
 INV_X1 _2783_ (.A(_2374_),
    .ZN(_1842_));
 NOR2_X2 _2784_ (.A1(net137),
    .A2(_1842_),
    .ZN(_1843_));
 NAND2_X1 _2785_ (.A1(_1645_),
    .A2(_1843_),
    .ZN(_1844_));
 MUX2_X1 _2786_ (.A(_1758_),
    .B(_1773_),
    .S(_1620_),
    .Z(_1845_));
 INV_X1 _2787_ (.A(_1845_),
    .ZN(_1846_));
 NAND2_X1 _2788_ (.A1(_1846_),
    .A2(net111),
    .ZN(_1847_));
 INV_X1 _2789_ (.A(_1784_),
    .ZN(_1848_));
 NAND2_X1 _2790_ (.A1(_1848_),
    .A2(_1546_),
    .ZN(_1849_));
 NAND2_X1 _2791_ (.A1(_1802_),
    .A2(net129),
    .ZN(_1850_));
 NAND3_X1 _2792_ (.A1(_1849_),
    .A2(_1576_),
    .A3(_1850_),
    .ZN(_1851_));
 NAND3_X1 _2793_ (.A1(_1847_),
    .A2(_1643_),
    .A3(_1851_),
    .ZN(_1852_));
 TAPCELL_X1 PHY_78 ();
 INV_X1 _2795_ (.A(net47),
    .ZN(_1854_));
 NOR2_X1 _2796_ (.A1(net123),
    .A2(_1854_),
    .ZN(_1855_));
 NAND2_X1 _2797_ (.A1(_1571_),
    .A2(_1855_),
    .ZN(_1856_));
 AND2_X1 _2798_ (.A1(net90),
    .A2(net46),
    .ZN(_1857_));
 NAND2_X1 _2799_ (.A1(_1571_),
    .A2(_1857_),
    .ZN(_1858_));
 MUX2_X1 _2800_ (.A(_1856_),
    .B(_1858_),
    .S(net93),
    .Z(_1859_));
 MUX2_X1 _2801_ (.A(_1822_),
    .B(_1859_),
    .S(_1546_),
    .Z(_1860_));
 MUX2_X1 _2802_ (.A(_1829_),
    .B(_1745_),
    .S(net145),
    .Z(_1861_));
 MUX2_X1 _2803_ (.A(_1860_),
    .B(_1861_),
    .S(_1576_),
    .Z(_1862_));
 AOI21_X1 _2804_ (.A(_1814_),
    .B1(_1862_),
    .B2(net89),
    .ZN(_1863_));
 NAND2_X1 _2805_ (.A1(_1852_),
    .A2(_1863_),
    .ZN(_1864_));
 NAND3_X1 _2806_ (.A1(_1627_),
    .A2(_1844_),
    .A3(_1864_),
    .ZN(_1865_));
 NAND2_X1 _2807_ (.A1(_1864_),
    .A2(_1844_),
    .ZN(_1866_));
 NAND2_X1 _2808_ (.A1(_1733_),
    .A2(_1866_),
    .ZN(_1867_));
 NAND2_X1 _2809_ (.A1(_1865_),
    .A2(_1867_),
    .ZN(_2012_));
 NAND2_X1 _2810_ (.A1(net101),
    .A2(net46),
    .ZN(_1868_));
 XNOR2_X2 _2811_ (.A(_1648_),
    .B(_1868_),
    .ZN(_2013_));
 NAND2_X1 _2812_ (.A1(_1830_),
    .A2(_1576_),
    .ZN(_1869_));
 INV_X1 _2813_ (.A(net45),
    .ZN(_1870_));
 NOR2_X1 _2814_ (.A1(net123),
    .A2(_1870_),
    .ZN(_1871_));
 INV_X1 _2815_ (.A(_1871_),
    .ZN(_1872_));
 OAI21_X1 _2816_ (.A(_1617_),
    .B1(_1570_),
    .B2(_1872_),
    .ZN(_1873_));
 INV_X1 _2817_ (.A(net44),
    .ZN(_1874_));
 NOR2_X1 _2818_ (.A1(net123),
    .A2(_1874_),
    .ZN(_1875_));
 INV_X1 _2819_ (.A(_1875_),
    .ZN(_1876_));
 NOR2_X1 _2820_ (.A1(_1570_),
    .A2(_1876_),
    .ZN(_1877_));
 OAI21_X1 _2821_ (.A(_1873_),
    .B1(_1877_),
    .B2(_1617_),
    .ZN(_1878_));
 OR2_X1 _2822_ (.A1(_1878_),
    .A2(net129),
    .ZN(_1879_));
 OAI21_X1 _2823_ (.A(_1879_),
    .B1(net102),
    .B2(_1859_),
    .ZN(_1880_));
 OAI21_X1 _2824_ (.A(_1869_),
    .B1(_1576_),
    .B2(_1880_),
    .ZN(_1881_));
 AOI21_X1 _2825_ (.A(_1814_),
    .B1(_1881_),
    .B2(net89),
    .ZN(_1882_));
 OAI21_X1 _2826_ (.A(_1882_),
    .B1(_1787_),
    .B2(net89),
    .ZN(_1883_));
 INV_X1 _2827_ (.A(_1843_),
    .ZN(_1884_));
 NOR2_X1 _2828_ (.A1(_1806_),
    .A2(_1643_),
    .ZN(_1885_));
 INV_X1 _2829_ (.A(_1885_),
    .ZN(_1886_));
 OAI21_X1 _2830_ (.A(_1883_),
    .B1(_1884_),
    .B2(_1886_),
    .ZN(_1887_));
 XNOR2_X1 _2831_ (.A(_1887_),
    .B(_1733_),
    .ZN(_2018_));
 NAND2_X1 _2832_ (.A1(net101),
    .A2(net44),
    .ZN(_1888_));
 XNOR2_X2 _2833_ (.A(_1648_),
    .B(_1888_),
    .ZN(_2017_));
 NAND2_X1 _2834_ (.A1(_1849_),
    .A2(_1850_),
    .ZN(_1889_));
 NAND2_X1 _2835_ (.A1(_1889_),
    .A2(net111),
    .ZN(_1890_));
 OAI21_X1 _2836_ (.A(_1890_),
    .B1(net105),
    .B2(_1637_),
    .ZN(_1891_));
 NOR2_X1 _2837_ (.A1(_1891_),
    .A2(_1643_),
    .ZN(_1892_));
 NAND2_X1 _2838_ (.A1(_1892_),
    .A2(_1843_),
    .ZN(_1893_));
 NAND2_X1 _2839_ (.A1(_1861_),
    .A2(net105),
    .ZN(_1894_));
 OAI21_X1 _2840_ (.A(_1894_),
    .B1(_1846_),
    .B2(net105),
    .ZN(_1895_));
 TAPCELL_X1 PHY_77 ();
 NAND2_X1 _2842_ (.A1(_1895_),
    .A2(_1643_),
    .ZN(_1897_));
 NAND2_X1 _2843_ (.A1(_1860_),
    .A2(_1576_),
    .ZN(_1898_));
 TAPCELL_X1 PHY_76 ();
 INV_X1 _2845_ (.A(net43),
    .ZN(_1900_));
 NOR2_X1 _2846_ (.A1(net109),
    .A2(_1900_),
    .ZN(_1901_));
 AND2_X1 _2847_ (.A1(_1571_),
    .A2(_1901_),
    .ZN(_1902_));
 NAND2_X1 _2848_ (.A1(_1902_),
    .A2(_1617_),
    .ZN(_1903_));
 NAND2_X1 _2849_ (.A1(net90),
    .A2(net42),
    .ZN(_1904_));
 INV_X1 _2850_ (.A(_1904_),
    .ZN(_1905_));
 NAND2_X1 _2851_ (.A1(_1571_),
    .A2(_1905_),
    .ZN(_1906_));
 OAI21_X1 _2852_ (.A(_1903_),
    .B1(_1617_),
    .B2(_1906_),
    .ZN(_1907_));
 NAND2_X1 _2853_ (.A1(_1907_),
    .A2(net103),
    .ZN(_1908_));
 OAI21_X1 _2854_ (.A(_1908_),
    .B1(net103),
    .B2(_1878_),
    .ZN(_1909_));
 OAI21_X1 _2855_ (.A(_1898_),
    .B1(_1576_),
    .B2(_1909_),
    .ZN(_1910_));
 AOI21_X1 _2856_ (.A(_1814_),
    .B1(_1910_),
    .B2(net89),
    .ZN(_1911_));
 NAND2_X1 _2857_ (.A1(_1897_),
    .A2(_1911_),
    .ZN(_1912_));
 NAND3_X1 _2858_ (.A1(_1627_),
    .A2(_1893_),
    .A3(_1912_),
    .ZN(_1913_));
 NAND2_X1 _2859_ (.A1(_1893_),
    .A2(_1912_),
    .ZN(_1914_));
 NAND2_X1 _2860_ (.A1(_1914_),
    .A2(_1733_),
    .ZN(_1915_));
 NAND2_X1 _2861_ (.A1(_1913_),
    .A2(_1915_),
    .ZN(_2022_));
 NAND2_X1 _2862_ (.A1(net101),
    .A2(net42),
    .ZN(_1916_));
 XNOR2_X2 _2863_ (.A(_1648_),
    .B(_1916_),
    .ZN(_2021_));
 NAND3_X1 _2864_ (.A1(_1836_),
    .A2(net89),
    .A3(_1843_),
    .ZN(_1917_));
 INV_X1 _2865_ (.A(net39),
    .ZN(_1918_));
 NOR2_X1 _2866_ (.A1(net123),
    .A2(_1918_),
    .ZN(_1919_));
 INV_X1 _2867_ (.A(_1919_),
    .ZN(_1920_));
 NOR2_X1 _2868_ (.A1(_1570_),
    .A2(_1920_),
    .ZN(_1921_));
 NAND2_X1 _2869_ (.A1(_1921_),
    .A2(_1617_),
    .ZN(_1922_));
 NAND2_X1 _2870_ (.A1(net90),
    .A2(net28),
    .ZN(_1923_));
 INV_X1 _2871_ (.A(_1923_),
    .ZN(_1924_));
 NAND2_X1 _2872_ (.A1(_1571_),
    .A2(_1924_),
    .ZN(_1925_));
 OAI21_X1 _2873_ (.A(_1922_),
    .B1(_1617_),
    .B2(_1925_),
    .ZN(_1926_));
 AOI21_X1 _2874_ (.A(_1576_),
    .B1(_1926_),
    .B2(net103),
    .ZN(_1927_));
 NAND2_X1 _2875_ (.A1(_1907_),
    .A2(net129),
    .ZN(_1928_));
 NAND2_X1 _2876_ (.A1(_1927_),
    .A2(_1928_),
    .ZN(_1929_));
 OAI21_X1 _2877_ (.A(_1929_),
    .B1(_1880_),
    .B2(net105),
    .ZN(_1930_));
 AOI21_X1 _2878_ (.A(_1814_),
    .B1(_1930_),
    .B2(net89),
    .ZN(_1931_));
 INV_X1 _2879_ (.A(_1832_),
    .ZN(_1932_));
 OAI21_X1 _2880_ (.A(_1931_),
    .B1(_1932_),
    .B2(net89),
    .ZN(_1933_));
 NAND3_X1 _2881_ (.A1(_1627_),
    .A2(_1917_),
    .A3(_1933_),
    .ZN(_1934_));
 NAND2_X1 _2882_ (.A1(_1917_),
    .A2(_1933_),
    .ZN(_1935_));
 NAND2_X1 _2883_ (.A1(_1935_),
    .A2(_1733_),
    .ZN(_1936_));
 NAND2_X1 _2884_ (.A1(_1934_),
    .A2(_1936_),
    .ZN(_2027_));
 NAND2_X1 _2885_ (.A1(net101),
    .A2(net28),
    .ZN(_0000_));
 XNOR2_X2 _2886_ (.A(_1648_),
    .B(_0000_),
    .ZN(_2026_));
 INV_X2 _2887_ (.A(_2362_),
    .ZN(_2370_));
 AOI21_X4 _2888_ (.A(_1575_),
    .B1(_2370_),
    .B2(_1553_),
    .ZN(_2373_));
 INV_X1 _2889_ (.A(_2353_),
    .ZN(_0001_));
 NAND2_X1 _2890_ (.A1(_2355_),
    .A2(_2031_),
    .ZN(_0002_));
 INV_X1 _2891_ (.A(_2354_),
    .ZN(_0003_));
 AOI21_X2 _2892_ (.A(_0001_),
    .B1(_0002_),
    .B2(_0003_),
    .ZN(_0004_));
 NOR2_X2 _2893_ (.A1(_2352_),
    .A2(_0004_),
    .ZN(_2028_));
 INV_X1 _2894_ (.A(_2336_),
    .ZN(_0005_));
 INV_X1 _2895_ (.A(_2337_),
    .ZN(_0006_));
 INV_X1 _2896_ (.A(_2340_),
    .ZN(_0007_));
 INV_X1 _2897_ (.A(_2344_),
    .ZN(_0008_));
 INV_X2 _2898_ (.A(_2345_),
    .ZN(_0009_));
 INV_X1 _2899_ (.A(_2348_),
    .ZN(_0010_));
 OAI21_X1 _2900_ (.A(_0008_),
    .B1(_0009_),
    .B2(_0010_),
    .ZN(_0011_));
 INV_X1 _2901_ (.A(_0011_),
    .ZN(_0012_));
 NAND2_X1 _2902_ (.A1(_2337_),
    .A2(_2341_),
    .ZN(_0013_));
 OAI221_X1 _2903_ (.A(_0005_),
    .B1(_0006_),
    .B2(_0007_),
    .C1(_0012_),
    .C2(_0013_),
    .ZN(_0014_));
 INV_X1 _2904_ (.A(_2028_),
    .ZN(_0015_));
 INV_X1 _2905_ (.A(_2349_),
    .ZN(_0016_));
 NOR3_X1 _2906_ (.A1(_0013_),
    .A2(_0009_),
    .A3(_0016_),
    .ZN(_0017_));
 AOI21_X2 _2907_ (.A(_0014_),
    .B1(_0015_),
    .B2(_0017_),
    .ZN(_2016_));
 INV_X1 _2908_ (.A(_2320_),
    .ZN(_0018_));
 INV_X1 _2909_ (.A(_2321_),
    .ZN(_0019_));
 INV_X1 _2910_ (.A(_2324_),
    .ZN(_0020_));
 INV_X1 _2911_ (.A(_2328_),
    .ZN(_0021_));
 INV_X1 _2912_ (.A(_2329_),
    .ZN(_0022_));
 INV_X1 _2913_ (.A(_2332_),
    .ZN(_0023_));
 OAI21_X1 _2914_ (.A(_0021_),
    .B1(_0022_),
    .B2(_0023_),
    .ZN(_0024_));
 INV_X1 _2915_ (.A(_0024_),
    .ZN(_0025_));
 NAND2_X1 _2916_ (.A1(_2321_),
    .A2(_2325_),
    .ZN(_0026_));
 OAI221_X1 _2917_ (.A(_0018_),
    .B1(_0019_),
    .B2(_0020_),
    .C1(_0025_),
    .C2(_0026_),
    .ZN(_0027_));
 INV_X2 _2918_ (.A(_2016_),
    .ZN(_0028_));
 NAND2_X1 _2919_ (.A1(_2329_),
    .A2(_2333_),
    .ZN(_0029_));
 NOR2_X1 _2920_ (.A1(_0026_),
    .A2(_0029_),
    .ZN(_0030_));
 AOI21_X4 _2921_ (.A(_0027_),
    .B1(_0028_),
    .B2(_0030_),
    .ZN(_2006_));
 NAND2_X1 _2922_ (.A1(_2313_),
    .A2(_2317_),
    .ZN(_0031_));
 OR2_X4 _2923_ (.A1(_0031_),
    .A2(_2006_),
    .ZN(_0032_));
 INV_X1 _2924_ (.A(_2312_),
    .ZN(_0033_));
 NAND2_X1 _2925_ (.A1(_2313_),
    .A2(_2316_),
    .ZN(_0034_));
 NAND3_X4 _2926_ (.A1(_0032_),
    .A2(_0033_),
    .A3(_0034_),
    .ZN(_2001_));
 NAND3_X4 _2927_ (.A1(_2001_),
    .A2(_2307_),
    .A3(_2309_),
    .ZN(_0035_));
 INV_X1 _2928_ (.A(_2306_),
    .ZN(_0036_));
 NAND2_X1 _2929_ (.A1(_2307_),
    .A2(_2308_),
    .ZN(_0037_));
 NAND3_X4 _2930_ (.A1(_0035_),
    .A2(_0036_),
    .A3(_0037_),
    .ZN(_0038_));
 INV_X4 _2931_ (.A(_0038_),
    .ZN(_1996_));
 INV_X1 _2932_ (.A(_2274_),
    .ZN(_0039_));
 INV_X1 _2933_ (.A(_2275_),
    .ZN(_0040_));
 INV_X1 _2934_ (.A(_2276_),
    .ZN(_0041_));
 OAI21_X1 _2935_ (.A(_0039_),
    .B1(_0040_),
    .B2(_0041_),
    .ZN(_0042_));
 INV_X1 _2936_ (.A(_2280_),
    .ZN(_0043_));
 INV_X1 _2937_ (.A(_2281_),
    .ZN(_0044_));
 INV_X1 _2938_ (.A(_2282_),
    .ZN(_0045_));
 INV_X1 _2939_ (.A(_2298_),
    .ZN(_0046_));
 INV_X1 _2940_ (.A(_2299_),
    .ZN(_0047_));
 INV_X1 _2941_ (.A(_2302_),
    .ZN(_0048_));
 OAI21_X1 _2942_ (.A(_0046_),
    .B1(_0047_),
    .B2(_0048_),
    .ZN(_0049_));
 INV_X1 _2943_ (.A(_0049_),
    .ZN(_0050_));
 NAND2_X1 _2944_ (.A1(_2299_),
    .A2(_2303_),
    .ZN(_0051_));
 OAI21_X4 _2945_ (.A(_0050_),
    .B1(_1996_),
    .B2(_0051_),
    .ZN(_1991_));
 NAND2_X1 _2946_ (.A1(_2293_),
    .A2(_2295_),
    .ZN(_0052_));
 INV_X1 _2947_ (.A(_0052_),
    .ZN(_0053_));
 NAND2_X4 _2948_ (.A1(_0053_),
    .A2(_1991_),
    .ZN(_0054_));
 INV_X1 _2949_ (.A(_2292_),
    .ZN(_0055_));
 NAND2_X1 _2950_ (.A1(_2293_),
    .A2(_2294_),
    .ZN(_0056_));
 NAND3_X4 _2951_ (.A1(_0054_),
    .A2(_0055_),
    .A3(_0056_),
    .ZN(_1986_));
 NAND2_X1 _2952_ (.A1(_2287_),
    .A2(_2289_),
    .ZN(_0057_));
 INV_X1 _2953_ (.A(_0057_),
    .ZN(_0058_));
 AND2_X4 _2954_ (.A1(_1986_),
    .A2(_0058_),
    .ZN(_0059_));
 INV_X1 _2955_ (.A(_2286_),
    .ZN(_0060_));
 INV_X1 _2956_ (.A(_2287_),
    .ZN(_0061_));
 INV_X1 _2957_ (.A(_2288_),
    .ZN(_0062_));
 OAI21_X1 _2958_ (.A(_0060_),
    .B1(_0061_),
    .B2(_0062_),
    .ZN(_0063_));
 NOR2_X4 _2959_ (.A1(_0063_),
    .A2(_0059_),
    .ZN(_0064_));
 NAND2_X1 _2960_ (.A1(_2281_),
    .A2(_2283_),
    .ZN(_0065_));
 OAI221_X2 _2961_ (.A(_0043_),
    .B1(_0044_),
    .B2(_0045_),
    .C1(_0064_),
    .C2(_0065_),
    .ZN(_1976_));
 NAND2_X1 _2962_ (.A1(_2275_),
    .A2(_2277_),
    .ZN(_0066_));
 INV_X1 _2963_ (.A(_0066_),
    .ZN(_0067_));
 AOI21_X2 _2964_ (.A(_0042_),
    .B1(_1976_),
    .B2(_0067_),
    .ZN(_1971_));
 INV_X1 _2965_ (.A(_0029_),
    .ZN(_0068_));
 AOI21_X1 _2966_ (.A(_0024_),
    .B1(_0028_),
    .B2(_0068_),
    .ZN(_2011_));
 NOR3_X1 _2967_ (.A1(_2028_),
    .A2(_0009_),
    .A3(_0016_),
    .ZN(_0069_));
 NOR2_X1 _2968_ (.A1(_0069_),
    .A2(_0011_),
    .ZN(_2023_));
 INV_X2 _2969_ (.A(_1980_),
    .ZN(_0070_));
 INV_X1 _2970_ (.A(_1979_),
    .ZN(_0071_));
 NAND2_X1 _2971_ (.A1(_0071_),
    .A2(_0040_),
    .ZN(_0072_));
 NAND2_X1 _2972_ (.A1(_1979_),
    .A2(_2275_),
    .ZN(_0073_));
 AOI21_X4 _2973_ (.A(_0070_),
    .B1(_0072_),
    .B2(_0073_),
    .ZN(_0074_));
 INV_X1 _2974_ (.A(_1974_),
    .ZN(_0075_));
 NAND3_X2 _2975_ (.A1(_1622_),
    .A2(_1623_),
    .A3(_0075_),
    .ZN(_0076_));
 TAPCELL_X1 PHY_75 ();
 NAND3_X4 _2977_ (.A1(_0074_),
    .A2(_0076_),
    .A3(_1975_),
    .ZN(_0078_));
 XNOR2_X2 _2978_ (.A(_0044_),
    .B(_1984_),
    .ZN(_0079_));
 INV_X1 _2979_ (.A(_1985_),
    .ZN(_0080_));
 NOR2_X1 _2980_ (.A1(_0079_),
    .A2(_0080_),
    .ZN(_0081_));
 XNOR2_X1 _2981_ (.A(_1989_),
    .B(_2287_),
    .ZN(_0082_));
 NAND2_X1 _2982_ (.A1(_0082_),
    .A2(_1990_),
    .ZN(_0083_));
 INV_X1 _2983_ (.A(_0083_),
    .ZN(_0084_));
 NAND2_X1 _2984_ (.A1(_0081_),
    .A2(_0084_),
    .ZN(_0085_));
 NOR2_X4 _2985_ (.A1(_0085_),
    .A2(_0078_),
    .ZN(_0086_));
 XNOR2_X1 _2986_ (.A(_2004_),
    .B(_2307_),
    .ZN(_0087_));
 INV_X1 _2987_ (.A(_0087_),
    .ZN(_0088_));
 INV_X1 _2988_ (.A(_2005_),
    .ZN(_0089_));
 NOR2_X1 _2989_ (.A1(_0088_),
    .A2(_0089_),
    .ZN(_0090_));
 INV_X1 _2990_ (.A(_2313_),
    .ZN(_0091_));
 NAND2_X1 _2991_ (.A1(_0091_),
    .A2(_2009_),
    .ZN(_0092_));
 INV_X1 _2992_ (.A(_2009_),
    .ZN(_0093_));
 NAND2_X1 _2993_ (.A1(_0093_),
    .A2(_2313_),
    .ZN(_0094_));
 NAND2_X2 _2994_ (.A1(_0092_),
    .A2(_0094_),
    .ZN(_0095_));
 NAND2_X1 _2995_ (.A1(_0095_),
    .A2(_2010_),
    .ZN(_0096_));
 INV_X1 _2996_ (.A(_0096_),
    .ZN(_0097_));
 NAND2_X1 _2997_ (.A1(_0090_),
    .A2(_0097_),
    .ZN(_0098_));
 INV_X1 _2998_ (.A(_1994_),
    .ZN(_0099_));
 NAND2_X1 _2999_ (.A1(_0099_),
    .A2(_2293_),
    .ZN(_0100_));
 INV_X1 _3000_ (.A(_2293_),
    .ZN(_0101_));
 NAND2_X1 _3001_ (.A1(_0101_),
    .A2(_1994_),
    .ZN(_0102_));
 TAPCELL_X1 PHY_74 ();
 NAND3_X1 _3003_ (.A1(_0100_),
    .A2(_0102_),
    .A3(_1995_),
    .ZN(_0104_));
 INV_X1 _3004_ (.A(_1999_),
    .ZN(_0105_));
 NAND2_X1 _3005_ (.A1(_0105_),
    .A2(_0047_),
    .ZN(_0106_));
 NAND2_X1 _3006_ (.A1(_1999_),
    .A2(_2299_),
    .ZN(_0107_));
 NAND3_X1 _3007_ (.A1(_0106_),
    .A2(_2000_),
    .A3(_0107_),
    .ZN(_0108_));
 NOR2_X1 _3008_ (.A1(_0104_),
    .A2(_0108_),
    .ZN(_0109_));
 INV_X1 _3009_ (.A(_0109_),
    .ZN(_0110_));
 NOR2_X1 _3010_ (.A1(_0098_),
    .A2(_0110_),
    .ZN(_0111_));
 NAND2_X4 _3011_ (.A1(_0086_),
    .A2(_0111_),
    .ZN(_0112_));
 INV_X1 _3012_ (.A(_2024_),
    .ZN(_0113_));
 NAND2_X1 _3013_ (.A1(_0113_),
    .A2(_2337_),
    .ZN(_0114_));
 NAND2_X1 _3014_ (.A1(_0006_),
    .A2(_2024_),
    .ZN(_0115_));
 NAND2_X2 _3015_ (.A1(_0114_),
    .A2(_0115_),
    .ZN(_0116_));
 NAND2_X1 _3016_ (.A1(_0116_),
    .A2(_2025_),
    .ZN(_0117_));
 INV_X1 _3017_ (.A(_2029_),
    .ZN(_0118_));
 NAND2_X1 _3018_ (.A1(_0118_),
    .A2(_2345_),
    .ZN(_0119_));
 NAND2_X1 _3019_ (.A1(_0009_),
    .A2(_2029_),
    .ZN(_0120_));
 NAND2_X2 _3020_ (.A1(_0119_),
    .A2(_0120_),
    .ZN(_0121_));
 NAND2_X1 _3021_ (.A1(_0121_),
    .A2(_2030_),
    .ZN(_0122_));
 NOR2_X1 _3022_ (.A1(_0117_),
    .A2(_0122_),
    .ZN(_0123_));
 INV_X1 _3023_ (.A(_2019_),
    .ZN(_0124_));
 NAND2_X1 _3024_ (.A1(_0124_),
    .A2(_2329_),
    .ZN(_0125_));
 NAND2_X1 _3025_ (.A1(_0022_),
    .A2(_2019_),
    .ZN(_0126_));
 NAND2_X1 _3026_ (.A1(_0125_),
    .A2(_0126_),
    .ZN(_0127_));
 NAND2_X1 _3027_ (.A1(_0127_),
    .A2(_2020_),
    .ZN(_0128_));
 INV_X1 _3028_ (.A(_2014_),
    .ZN(_0129_));
 NAND2_X1 _3029_ (.A1(_0129_),
    .A2(_0019_),
    .ZN(_0130_));
 TAPCELL_X1 PHY_73 ();
 NAND2_X1 _3031_ (.A1(_2014_),
    .A2(_2321_),
    .ZN(_0132_));
 NAND3_X1 _3032_ (.A1(_0130_),
    .A2(_2015_),
    .A3(_0132_),
    .ZN(_0133_));
 NOR2_X2 _3033_ (.A1(_0128_),
    .A2(_0133_),
    .ZN(_0134_));
 NAND2_X1 _3034_ (.A1(_0123_),
    .A2(_0134_),
    .ZN(_0135_));
 XNOR2_X2 _3035_ (.A(_2034_),
    .B(_2353_),
    .ZN(_0136_));
 TAPCELL_X1 PHY_72 ();
 INV_X1 _3037_ (.A(_2035_),
    .ZN(_0138_));
 NAND2_X1 _3038_ (.A1(_0136_),
    .A2(_0138_),
    .ZN(_0139_));
 INV_X1 _3039_ (.A(_2038_),
    .ZN(_0140_));
 INV_X1 _3040_ (.A(_2041_),
    .ZN(_0141_));
 NAND2_X1 _3041_ (.A1(_0140_),
    .A2(_0141_),
    .ZN(_0142_));
 OR2_X1 _3042_ (.A1(_0139_),
    .A2(_0142_),
    .ZN(_0143_));
 NOR2_X1 _3043_ (.A1(_0135_),
    .A2(_0143_),
    .ZN(_0144_));
 NOR2_X4 _3044_ (.A1(_0144_),
    .A2(_0112_),
    .ZN(_2068_));
 NAND3_X1 _3045_ (.A1(_0125_),
    .A2(_0126_),
    .A3(_2015_),
    .ZN(_0145_));
 AND2_X1 _3046_ (.A1(_0130_),
    .A2(_0132_),
    .ZN(_0146_));
 NAND2_X1 _3047_ (.A1(_0145_),
    .A2(_0146_),
    .ZN(_0147_));
 INV_X1 _3048_ (.A(_2025_),
    .ZN(_0148_));
 OAI21_X1 _3049_ (.A(_0116_),
    .B1(_0121_),
    .B2(_0148_),
    .ZN(_0149_));
 AOI21_X1 _3050_ (.A(_0147_),
    .B1(_0134_),
    .B2(_0149_),
    .ZN(_0150_));
 OAI21_X1 _3051_ (.A(_0136_),
    .B1(_0140_),
    .B2(_2035_),
    .ZN(_0151_));
 NAND3_X1 _3052_ (.A1(_0123_),
    .A2(_0134_),
    .A3(_0151_),
    .ZN(_0152_));
 NAND2_X1 _3053_ (.A1(_0150_),
    .A2(_0152_),
    .ZN(_0153_));
 INV_X1 _3054_ (.A(_0153_),
    .ZN(_0154_));
 NAND2_X2 _3055_ (.A1(_2068_),
    .A2(_0154_),
    .ZN(_0155_));
 OAI21_X1 _3056_ (.A(_0087_),
    .B1(_0095_),
    .B2(_0089_),
    .ZN(_0156_));
 NAND2_X1 _3057_ (.A1(_0109_),
    .A2(_0156_),
    .ZN(_0157_));
 NAND2_X2 _3058_ (.A1(_0100_),
    .A2(_0102_),
    .ZN(_0158_));
 INV_X1 _3059_ (.A(_0158_),
    .ZN(_0159_));
 AND2_X1 _3060_ (.A1(_0106_),
    .A2(_0107_),
    .ZN(_0160_));
 INV_X1 _3061_ (.A(_1995_),
    .ZN(_0161_));
 OAI21_X1 _3062_ (.A(_0159_),
    .B1(_0160_),
    .B2(_0161_),
    .ZN(_0162_));
 INV_X1 _3063_ (.A(_0162_),
    .ZN(_0163_));
 NAND2_X1 _3064_ (.A1(_0157_),
    .A2(_0163_),
    .ZN(_0164_));
 NAND2_X1 _3065_ (.A1(_0164_),
    .A2(_0086_),
    .ZN(_0165_));
 NAND2_X1 _3066_ (.A1(_0072_),
    .A2(_0073_),
    .ZN(_0166_));
 INV_X1 _3067_ (.A(_0166_),
    .ZN(_0167_));
 NAND2_X1 _3068_ (.A1(_0167_),
    .A2(_1975_),
    .ZN(_0168_));
 NAND2_X1 _3069_ (.A1(_0168_),
    .A2(_0076_),
    .ZN(_0169_));
 NAND2_X2 _3070_ (.A1(_1975_),
    .A2(_0076_),
    .ZN(_0170_));
 INV_X4 _3071_ (.A(_0074_),
    .ZN(_0171_));
 NOR2_X4 _3072_ (.A1(_0171_),
    .A2(_0170_),
    .ZN(_0172_));
 INV_X1 _3073_ (.A(_0079_),
    .ZN(_0173_));
 OAI21_X1 _3074_ (.A(_0173_),
    .B1(_0082_),
    .B2(_0080_),
    .ZN(_0174_));
 AOI21_X1 _3075_ (.A(_0169_),
    .B1(_0172_),
    .B2(_0174_),
    .ZN(_0175_));
 NAND3_X1 _3076_ (.A1(_0165_),
    .A2(_0175_),
    .A3(_0112_),
    .ZN(_0176_));
 NAND2_X2 _3077_ (.A1(_0155_),
    .A2(_0176_),
    .ZN(_0177_));
 INV_X2 _3078_ (.A(_0177_),
    .ZN(_2093_));
 INV_X1 _3079_ (.A(net32),
    .ZN(_2267_));
 INV_X1 _3080_ (.A(net33),
    .ZN(_1941_));
 NOR2_X1 _3081_ (.A1(net118),
    .A2(_1941_),
    .ZN(_0178_));
 INV_X1 _3082_ (.A(_1938_),
    .ZN(_1942_));
 AOI21_X2 _3083_ (.A(_0178_),
    .B1(_1942_),
    .B2(net113),
    .ZN(_2088_));
 INV_X1 _3084_ (.A(net34),
    .ZN(_1949_));
 NAND2_X1 _3085_ (.A1(_1946_),
    .A2(net118),
    .ZN(_0179_));
 OAI21_X2 _3086_ (.A(_0179_),
    .B1(net34),
    .B2(_1542_),
    .ZN(_2084_));
 INV_X1 _3087_ (.A(net35),
    .ZN(_2211_));
 INV_X2 _3088_ (.A(_2215_),
    .ZN(_2212_));
 NAND2_X1 _3089_ (.A1(_2212_),
    .A2(net118),
    .ZN(_0180_));
 OAI21_X2 _3090_ (.A(_0180_),
    .B1(_2211_),
    .B2(net118),
    .ZN(_2073_));
 INV_X1 _3091_ (.A(_2073_),
    .ZN(_2077_));
 INV_X1 _3092_ (.A(net36),
    .ZN(_1953_));
 NAND2_X1 _3093_ (.A1(net90),
    .A2(_1958_),
    .ZN(_0181_));
 NAND2_X1 _3094_ (.A1(net101),
    .A2(_1953_),
    .ZN(_0182_));
 NAND2_X1 _3095_ (.A1(_0181_),
    .A2(_0182_),
    .ZN(_2069_));
 INV_X1 _3096_ (.A(_1962_),
    .ZN(_1967_));
 NAND2_X1 _3097_ (.A1(_1962_),
    .A2(net90),
    .ZN(_0183_));
 INV_X1 _3098_ (.A(net37),
    .ZN(_2202_));
 NAND2_X1 _3099_ (.A1(net101),
    .A2(_2202_),
    .ZN(_0184_));
 NAND2_X2 _3100_ (.A1(_0183_),
    .A2(_0184_),
    .ZN(_2139_));
 INV_X1 _3101_ (.A(_2139_),
    .ZN(_2060_));
 INV_X1 _3102_ (.A(net38),
    .ZN(_1966_));
 OAI21_X2 _3103_ (.A(_0183_),
    .B1(net38),
    .B2(net90),
    .ZN(_2059_));
 NAND2_X1 _3104_ (.A1(net90),
    .A2(_2195_),
    .ZN(_0185_));
 INV_X1 _3105_ (.A(net40),
    .ZN(_0186_));
 NAND2_X1 _3106_ (.A1(net101),
    .A2(_0186_),
    .ZN(_0187_));
 NAND2_X2 _3107_ (.A1(_0185_),
    .A2(_0187_),
    .ZN(_2142_));
 INV_X1 _3108_ (.A(_2142_),
    .ZN(_2145_));
 NAND2_X1 _3109_ (.A1(_0086_),
    .A2(_0110_),
    .ZN(_0188_));
 NAND3_X2 _3110_ (.A1(_0112_),
    .A2(_0188_),
    .A3(_0172_),
    .ZN(_0189_));
 INV_X4 _3111_ (.A(_2068_),
    .ZN(_2064_));
 INV_X1 _3112_ (.A(_0135_),
    .ZN(_0190_));
 NAND2_X1 _3113_ (.A1(_0190_),
    .A2(_0143_),
    .ZN(_0191_));
 NAND2_X1 _3114_ (.A1(_0191_),
    .A2(_0134_),
    .ZN(_0192_));
 OAI21_X4 _3115_ (.A(_0189_),
    .B1(_2064_),
    .B2(_0192_),
    .ZN(_2083_));
 INV_X1 _3116_ (.A(_2067_),
    .ZN(_2055_));
 INV_X1 _3117_ (.A(_0085_),
    .ZN(_0193_));
 NAND2_X4 _3118_ (.A1(_0193_),
    .A2(_0172_),
    .ZN(_0194_));
 AOI21_X2 _3119_ (.A(_0194_),
    .B1(_0191_),
    .B2(_0111_),
    .ZN(_2076_));
 NAND2_X1 _3120_ (.A1(_0190_),
    .A2(_0139_),
    .ZN(_0195_));
 AOI21_X1 _3121_ (.A(_0133_),
    .B1(_0134_),
    .B2(_0117_),
    .ZN(_0196_));
 NAND2_X1 _3122_ (.A1(_0195_),
    .A2(_0196_),
    .ZN(_0197_));
 NAND3_X1 _3123_ (.A1(_0109_),
    .A2(_0090_),
    .A3(_0097_),
    .ZN(_0198_));
 NOR2_X4 _3124_ (.A1(_0198_),
    .A2(_0194_),
    .ZN(_0199_));
 NAND2_X1 _3125_ (.A1(_0197_),
    .A2(_0199_),
    .ZN(_0200_));
 NOR2_X1 _3126_ (.A1(_0078_),
    .A2(_0081_),
    .ZN(_0201_));
 NOR2_X1 _3127_ (.A1(_0201_),
    .A2(_0170_),
    .ZN(_0202_));
 INV_X1 _3128_ (.A(_0104_),
    .ZN(_0203_));
 OAI21_X1 _3129_ (.A(_0203_),
    .B1(_0090_),
    .B2(_0108_),
    .ZN(_0204_));
 NAND2_X1 _3130_ (.A1(_0086_),
    .A2(_0204_),
    .ZN(_0205_));
 NAND2_X1 _3131_ (.A1(_0202_),
    .A2(_0205_),
    .ZN(_0206_));
 INV_X1 _3132_ (.A(_0206_),
    .ZN(_0207_));
 NAND2_X2 _3133_ (.A1(_0200_),
    .A2(_0207_),
    .ZN(_0208_));
 NAND2_X4 _3134_ (.A1(_0144_),
    .A2(_0199_),
    .ZN(_0209_));
 INV_X4 _3135_ (.A(_0209_),
    .ZN(_0210_));
 NOR2_X4 _3136_ (.A1(_0208_),
    .A2(_0210_),
    .ZN(_2087_));
 INV_X2 _3137_ (.A(_2083_),
    .ZN(_2080_));
 INV_X1 _3138_ (.A(_2143_),
    .ZN(_0211_));
 INV_X1 _3139_ (.A(_2094_),
    .ZN(_0212_));
 OAI21_X1 _3140_ (.A(_2090_),
    .B1(_0212_),
    .B2(_2095_),
    .ZN(_0213_));
 INV_X1 _3141_ (.A(_2089_),
    .ZN(_0214_));
 NAND2_X1 _3142_ (.A1(_0213_),
    .A2(_0214_),
    .ZN(_0215_));
 NAND2_X1 _3143_ (.A1(_2075_),
    .A2(_2051_),
    .ZN(_0216_));
 INV_X1 _3144_ (.A(_0216_),
    .ZN(_0217_));
 NAND2_X1 _3145_ (.A1(_0215_),
    .A2(_0217_),
    .ZN(_0218_));
 NAND2_X1 _3146_ (.A1(_2075_),
    .A2(_2085_),
    .ZN(_0219_));
 INV_X1 _3147_ (.A(_2078_),
    .ZN(_0220_));
 NAND2_X1 _3148_ (.A1(_0219_),
    .A2(_0220_),
    .ZN(_0221_));
 INV_X1 _3149_ (.A(_0221_),
    .ZN(_0222_));
 NAND2_X1 _3150_ (.A1(_0222_),
    .A2(_0218_),
    .ZN(_0223_));
 NAND2_X2 _3151_ (.A1(_0223_),
    .A2(_2067_),
    .ZN(_0224_));
 INV_X1 _3152_ (.A(_2070_),
    .ZN(_0225_));
 AOI21_X4 _3153_ (.A(_0211_),
    .B1(_0224_),
    .B2(_0225_),
    .ZN(_0226_));
 NAND2_X4 _3154_ (.A1(_0226_),
    .A2(_2139_),
    .ZN(_0227_));
 NAND2_X4 _3155_ (.A1(_0209_),
    .A2(_0227_),
    .ZN(_0228_));
 INV_X16 _3156_ (.A(_0228_),
    .ZN(_0229_));
 NAND2_X4 _3157_ (.A1(_2083_),
    .A2(_0229_),
    .ZN(_0230_));
 NAND2_X4 _3158_ (.A1(_0228_),
    .A2(_2098_),
    .ZN(_0231_));
 AND2_X4 _3159_ (.A1(_0231_),
    .A2(_0230_),
    .ZN(_0232_));
 TAPCELL_X1 PHY_71 ();
 TAPCELL_X1 PHY_70 ();
 INV_X1 _3162_ (.A(_2084_),
    .ZN(_2081_));
 AND3_X1 _3163_ (.A1(_2073_),
    .A2(_2096_),
    .A3(_2081_),
    .ZN(_2103_));
 INV_X1 _3164_ (.A(_2069_),
    .ZN(_2065_));
 NAND3_X1 _3165_ (.A1(_2103_),
    .A2(_2065_),
    .A3(_2060_),
    .ZN(_0234_));
 INV_X1 _3166_ (.A(_0234_),
    .ZN(_2099_));
 NAND3_X1 _3167_ (.A1(_2099_),
    .A2(_2146_),
    .A3(_0228_),
    .ZN(_2126_));
 INV_X1 _3168_ (.A(_2126_),
    .ZN(_2130_));
 TAPCELL_X1 PHY_69 ();
 TAPCELL_X1 PHY_68 ();
 NAND2_X1 _3171_ (.A1(net150),
    .A2(_2064_),
    .ZN(_0237_));
 OAI21_X1 _3172_ (.A(_0237_),
    .B1(_2105_),
    .B2(net150),
    .ZN(_2118_));
 XNOR2_X1 _3173_ (.A(_2060_),
    .B(_2104_),
    .ZN(_0238_));
 NOR2_X1 _3174_ (.A1(_0238_),
    .A2(_0229_),
    .ZN(_0239_));
 INV_X1 _3175_ (.A(_2116_),
    .ZN(_0240_));
 OAI21_X2 _3176_ (.A(_0239_),
    .B1(_0240_),
    .B2(_2105_),
    .ZN(_0241_));
 INV_X1 _3177_ (.A(_2102_),
    .ZN(_0242_));
 INV_X1 _3178_ (.A(_2101_),
    .ZN(_0243_));
 XNOR2_X1 _3179_ (.A(_2142_),
    .B(_0243_),
    .ZN(_0244_));
 INV_X1 _3180_ (.A(_0244_),
    .ZN(_0245_));
 NAND2_X1 _3181_ (.A1(_0245_),
    .A2(_0228_),
    .ZN(_0246_));
 NOR4_X2 _3182_ (.A1(_0241_),
    .A2(_0242_),
    .A3(_0229_),
    .A4(_0246_),
    .ZN(_2129_));
 XOR2_X2 _3183_ (.A(_0239_),
    .B(_2119_),
    .Z(_0247_));
 TAPCELL_X1 PHY_67 ();
 NAND2_X1 _3185_ (.A1(net150),
    .A2(_0177_),
    .ZN(_0249_));
 NAND2_X1 _3186_ (.A1(_0228_),
    .A2(_2108_),
    .ZN(_0250_));
 NAND2_X4 _3187_ (.A1(_0249_),
    .A2(_0250_),
    .ZN(_0251_));
 TAPCELL_X1 PHY_66 ();
 TAPCELL_X1 PHY_65 ();
 NAND2_X1 _3190_ (.A1(_0079_),
    .A2(net99),
    .ZN(_0254_));
 INV_X1 _3191_ (.A(_0254_),
    .ZN(_0255_));
 NAND2_X1 _3192_ (.A1(_0251_),
    .A2(_0255_),
    .ZN(_0256_));
 NAND2_X1 _3193_ (.A1(_0165_),
    .A2(_0175_),
    .ZN(_0257_));
 INV_X1 _3194_ (.A(_0257_),
    .ZN(_0258_));
 NAND2_X1 _3195_ (.A1(_0153_),
    .A2(_0199_),
    .ZN(_0259_));
 NAND2_X1 _3196_ (.A1(_0258_),
    .A2(_0259_),
    .ZN(_0260_));
 NAND3_X4 _3197_ (.A1(_0260_),
    .A2(_0209_),
    .A3(_0227_),
    .ZN(_0261_));
 INV_X1 _3198_ (.A(_2108_),
    .ZN(_0262_));
 NAND2_X4 _3199_ (.A1(_0228_),
    .A2(_0262_),
    .ZN(_0263_));
 NAND2_X4 _3200_ (.A1(_0261_),
    .A2(_0263_),
    .ZN(_0264_));
 TAPCELL_X1 PHY_64 ();
 TAPCELL_X1 PHY_63 ();
 INV_X4 _3203_ (.A(_2127_),
    .ZN(_0267_));
 TAPCELL_X1 PHY_62 ();
 NOR2_X1 _3205_ (.A1(net120),
    .A2(_1980_),
    .ZN(_0269_));
 NAND2_X1 _3206_ (.A1(_0264_),
    .A2(_0269_),
    .ZN(_0270_));
 NAND3_X1 _3207_ (.A1(_0208_),
    .A2(_0209_),
    .A3(_0227_),
    .ZN(_0271_));
 INV_X1 _3208_ (.A(_2110_),
    .ZN(_0272_));
 NAND2_X1 _3209_ (.A1(_0228_),
    .A2(_0272_),
    .ZN(_0273_));
 NAND2_X4 _3210_ (.A1(_0271_),
    .A2(_0273_),
    .ZN(_0274_));
 TAPCELL_X1 PHY_61 ();
 NAND3_X1 _3212_ (.A1(_0256_),
    .A2(_0270_),
    .A3(_0274_),
    .ZN(_0276_));
 TAPCELL_X1 PHY_60 ();
 XNOR2_X1 _3214_ (.A(_0061_),
    .B(_1989_),
    .ZN(_0278_));
 NAND2_X1 _3215_ (.A1(_0278_),
    .A2(net99),
    .ZN(_0279_));
 INV_X1 _3216_ (.A(_0279_),
    .ZN(_0280_));
 NAND2_X1 _3217_ (.A1(_0251_),
    .A2(_0280_),
    .ZN(_0281_));
 NOR2_X1 _3218_ (.A1(net120),
    .A2(_1985_),
    .ZN(_0282_));
 NAND2_X1 _3219_ (.A1(_0264_),
    .A2(_0282_),
    .ZN(_0283_));
 INV_X8 _3220_ (.A(_0274_),
    .ZN(_0284_));
 TAPCELL_X1 PHY_59 ();
 NAND3_X1 _3222_ (.A1(_0281_),
    .A2(_0283_),
    .A3(_0284_),
    .ZN(_0286_));
 NAND3_X1 _3223_ (.A1(_0276_),
    .A2(_0286_),
    .A3(net117),
    .ZN(_0287_));
 NAND2_X1 _3224_ (.A1(_0167_),
    .A2(_2127_),
    .ZN(_0288_));
 INV_X1 _3225_ (.A(_0288_),
    .ZN(_0289_));
 NAND2_X1 _3226_ (.A1(_0251_),
    .A2(_0289_),
    .ZN(_0290_));
 TAPCELL_X1 PHY_58 ();
 NOR2_X1 _3228_ (.A1(net120),
    .A2(_1975_),
    .ZN(_0292_));
 NAND2_X1 _3229_ (.A1(_0264_),
    .A2(_0292_),
    .ZN(_0293_));
 NAND3_X1 _3230_ (.A1(_0290_),
    .A2(_0293_),
    .A3(_0284_),
    .ZN(_0294_));
 INV_X8 _3231_ (.A(net114),
    .ZN(_0295_));
 TAPCELL_X1 PHY_57 ();
 TAPCELL_X1 PHY_56 ();
 NOR2_X1 _3234_ (.A1(_0076_),
    .A2(net120),
    .ZN(_0298_));
 INV_X1 _3235_ (.A(_0298_),
    .ZN(_0299_));
 OAI21_X1 _3236_ (.A(_0274_),
    .B1(_0264_),
    .B2(_0299_),
    .ZN(_0300_));
 NAND3_X1 _3237_ (.A1(_0294_),
    .A2(_0295_),
    .A3(_0300_),
    .ZN(_0301_));
 NAND2_X1 _3238_ (.A1(_0287_),
    .A2(_0301_),
    .ZN(_0302_));
 INV_X1 _3239_ (.A(_0302_),
    .ZN(_0303_));
 TAPCELL_X1 PHY_55 ();
 INV_X8 _3241_ (.A(net85),
    .ZN(_0305_));
 TAPCELL_X1 PHY_54 ();
 NOR2_X1 _3243_ (.A1(_0303_),
    .A2(_0305_),
    .ZN(_0307_));
 INV_X1 _3244_ (.A(_0307_),
    .ZN(_0308_));
 TAPCELL_X1 PHY_53 ();
 TAPCELL_X1 PHY_52 ();
 OAI21_X1 _3247_ (.A(_0247_),
    .B1(_0308_),
    .B2(_2120_),
    .ZN(_0311_));
 INV_X1 _3248_ (.A(_2123_),
    .ZN(_0312_));
 NAND2_X1 _3249_ (.A1(_0246_),
    .A2(_0312_),
    .ZN(_0313_));
 NAND3_X1 _3250_ (.A1(_0245_),
    .A2(_2123_),
    .A3(_0228_),
    .ZN(_0314_));
 NAND2_X4 _3251_ (.A1(_0313_),
    .A2(_0314_),
    .ZN(_0315_));
 INV_X1 _3252_ (.A(_2124_),
    .ZN(_0316_));
 NAND2_X4 _3253_ (.A1(_0315_),
    .A2(_0316_),
    .ZN(_0317_));
 NAND2_X1 _3254_ (.A1(_2038_),
    .A2(net99),
    .ZN(_0318_));
 NAND2_X1 _3255_ (.A1(_0251_),
    .A2(_0318_),
    .ZN(_0319_));
 NAND2_X1 _3256_ (.A1(_2035_),
    .A2(net99),
    .ZN(_0320_));
 NAND2_X1 _3257_ (.A1(_0264_),
    .A2(_0320_),
    .ZN(_0321_));
 TAPCELL_X1 PHY_51 ();
 NAND3_X1 _3259_ (.A1(_0319_),
    .A2(_0321_),
    .A3(_0284_),
    .ZN(_0323_));
 OR2_X1 _3260_ (.A1(_0136_),
    .A2(_0267_),
    .ZN(_0324_));
 NAND2_X1 _3261_ (.A1(_0251_),
    .A2(_0324_),
    .ZN(_0325_));
 NOR2_X1 _3262_ (.A1(_0267_),
    .A2(_2030_),
    .ZN(_0326_));
 INV_X1 _3263_ (.A(_0326_),
    .ZN(_0327_));
 NAND2_X1 _3264_ (.A1(_0264_),
    .A2(_0327_),
    .ZN(_0328_));
 TAPCELL_X1 PHY_50 ();
 NAND3_X1 _3266_ (.A1(_0325_),
    .A2(_0328_),
    .A3(_0274_),
    .ZN(_0330_));
 NAND3_X1 _3267_ (.A1(_0323_),
    .A2(_0330_),
    .A3(_0295_),
    .ZN(_0331_));
 NAND2_X1 _3268_ (.A1(_2041_),
    .A2(net100),
    .ZN(_0332_));
 INV_X1 _3269_ (.A(_0332_),
    .ZN(_0333_));
 NAND3_X1 _3270_ (.A1(_0274_),
    .A2(_0264_),
    .A3(_0333_),
    .ZN(_0334_));
 TAPCELL_X1 PHY_49 ();
 NAND2_X1 _3272_ (.A1(_0334_),
    .A2(net104),
    .ZN(_0336_));
 AND2_X1 _3273_ (.A1(_0331_),
    .A2(_0336_),
    .ZN(_0337_));
 TAPCELL_X1 PHY_48 ();
 TAPCELL_X1 PHY_47 ();
 NAND2_X1 _3276_ (.A1(_0337_),
    .A2(_0305_),
    .ZN(_0340_));
 NOR2_X2 _3277_ (.A1(net81),
    .A2(net83),
    .ZN(_0341_));
 AOI21_X1 _3278_ (.A(_0317_),
    .B1(_0340_),
    .B2(_0341_),
    .ZN(_0342_));
 NAND2_X1 _3279_ (.A1(_0311_),
    .A2(_0342_),
    .ZN(_0343_));
 INV_X8 _3280_ (.A(net82),
    .ZN(_0344_));
 TAPCELL_X1 PHY_46 ();
 NAND2_X1 _3282_ (.A1(_0158_),
    .A2(net99),
    .ZN(_0346_));
 NAND2_X1 _3283_ (.A1(_0251_),
    .A2(_0346_),
    .ZN(_0347_));
 NOR2_X1 _3284_ (.A1(_0267_),
    .A2(_1990_),
    .ZN(_0348_));
 INV_X1 _3285_ (.A(_0348_),
    .ZN(_0349_));
 NAND2_X1 _3286_ (.A1(_0264_),
    .A2(_0349_),
    .ZN(_0350_));
 NAND2_X1 _3287_ (.A1(_0347_),
    .A2(_0350_),
    .ZN(_0351_));
 NAND2_X1 _3288_ (.A1(_0351_),
    .A2(_0274_),
    .ZN(_0352_));
 TAPCELL_X1 PHY_45 ();
 NOR2_X1 _3290_ (.A1(_0160_),
    .A2(_0267_),
    .ZN(_0354_));
 NAND2_X1 _3291_ (.A1(_0251_),
    .A2(_0354_),
    .ZN(_0355_));
 NOR2_X2 _3292_ (.A1(net132),
    .A2(_1995_),
    .ZN(_0356_));
 NAND2_X1 _3293_ (.A1(_0264_),
    .A2(_0356_),
    .ZN(_0357_));
 NAND3_X1 _3294_ (.A1(_0355_),
    .A2(_0357_),
    .A3(_0284_),
    .ZN(_0358_));
 NAND2_X1 _3295_ (.A1(_0352_),
    .A2(_0358_),
    .ZN(_0359_));
 INV_X1 _3296_ (.A(_0359_),
    .ZN(_0360_));
 NAND2_X1 _3297_ (.A1(_0360_),
    .A2(_0295_),
    .ZN(_0361_));
 NAND2_X1 _3298_ (.A1(_0088_),
    .A2(net99),
    .ZN(_0362_));
 NAND2_X1 _3299_ (.A1(_0251_),
    .A2(_0362_),
    .ZN(_0363_));
 TAPCELL_X1 PHY_44 ();
 NOR2_X2 _3301_ (.A1(net120),
    .A2(_2000_),
    .ZN(_0365_));
 INV_X1 _3302_ (.A(_0365_),
    .ZN(_0366_));
 NAND2_X1 _3303_ (.A1(_0264_),
    .A2(_0366_),
    .ZN(_0367_));
 NAND2_X1 _3304_ (.A1(_0363_),
    .A2(_0367_),
    .ZN(_0368_));
 NAND2_X1 _3305_ (.A1(_0368_),
    .A2(_0274_),
    .ZN(_0369_));
 NOR2_X2 _3306_ (.A1(net120),
    .A2(_2005_),
    .ZN(_0370_));
 INV_X1 _3307_ (.A(_0370_),
    .ZN(_0371_));
 NAND2_X1 _3308_ (.A1(_0264_),
    .A2(_0371_),
    .ZN(_0372_));
 NOR2_X2 _3309_ (.A1(_0095_),
    .A2(net120),
    .ZN(_0373_));
 INV_X1 _3310_ (.A(_0373_),
    .ZN(_0374_));
 NAND3_X1 _3311_ (.A1(_0261_),
    .A2(_0263_),
    .A3(_0374_),
    .ZN(_0375_));
 NAND2_X1 _3312_ (.A1(_0372_),
    .A2(_0375_),
    .ZN(_0376_));
 NAND2_X1 _3313_ (.A1(_0376_),
    .A2(_0284_),
    .ZN(_0377_));
 NAND3_X1 _3314_ (.A1(_0369_),
    .A2(_0377_),
    .A3(net117),
    .ZN(_0378_));
 NAND2_X1 _3315_ (.A1(_0361_),
    .A2(_0378_),
    .ZN(_0379_));
 INV_X1 _3316_ (.A(_0379_),
    .ZN(_0380_));
 TAPCELL_X1 PHY_43 ();
 NAND2_X1 _3318_ (.A1(_0380_),
    .A2(_0305_),
    .ZN(_0382_));
 NOR2_X2 _3319_ (.A1(net120),
    .A2(_2010_),
    .ZN(_0383_));
 INV_X1 _3320_ (.A(_0383_),
    .ZN(_0384_));
 NAND2_X1 _3321_ (.A1(_0384_),
    .A2(_0264_),
    .ZN(_0385_));
 NOR2_X2 _3322_ (.A1(_0146_),
    .A2(net132),
    .ZN(_0386_));
 INV_X1 _3323_ (.A(_0386_),
    .ZN(_0387_));
 NAND3_X1 _3324_ (.A1(_0261_),
    .A2(_0263_),
    .A3(_0387_),
    .ZN(_0388_));
 NAND3_X1 _3325_ (.A1(_0385_),
    .A2(_0388_),
    .A3(_0274_),
    .ZN(_0389_));
 TAPCELL_X1 PHY_42 ();
 NOR2_X1 _3327_ (.A1(_0127_),
    .A2(_0267_),
    .ZN(_0391_));
 INV_X1 _3328_ (.A(_0391_),
    .ZN(_0392_));
 NAND2_X1 _3329_ (.A1(_0251_),
    .A2(_0392_),
    .ZN(_0393_));
 NOR2_X2 _3330_ (.A1(net132),
    .A2(_2015_),
    .ZN(_0394_));
 INV_X1 _3331_ (.A(_0394_),
    .ZN(_0395_));
 NAND2_X1 _3332_ (.A1(_0264_),
    .A2(_0395_),
    .ZN(_0396_));
 NAND2_X1 _3333_ (.A1(_0393_),
    .A2(_0396_),
    .ZN(_0397_));
 OAI21_X2 _3334_ (.A(_0389_),
    .B1(_0274_),
    .B2(_0397_),
    .ZN(_0398_));
 TAPCELL_X1 PHY_41 ();
 NAND2_X1 _3336_ (.A1(_0398_),
    .A2(_0295_),
    .ZN(_0400_));
 NOR2_X2 _3337_ (.A1(_0116_),
    .A2(net120),
    .ZN(_0401_));
 INV_X1 _3338_ (.A(_0401_),
    .ZN(_0402_));
 NAND2_X1 _3339_ (.A1(_0251_),
    .A2(_0402_),
    .ZN(_0403_));
 NOR2_X2 _3340_ (.A1(net132),
    .A2(_2020_),
    .ZN(_0404_));
 INV_X1 _3341_ (.A(_0404_),
    .ZN(_0405_));
 NAND2_X1 _3342_ (.A1(_0264_),
    .A2(_0405_),
    .ZN(_0406_));
 NAND2_X2 _3343_ (.A1(_0403_),
    .A2(_0406_),
    .ZN(_0407_));
 NAND2_X2 _3344_ (.A1(_0407_),
    .A2(_0274_),
    .ZN(_0408_));
 NOR2_X2 _3345_ (.A1(net132),
    .A2(_2025_),
    .ZN(_0409_));
 INV_X1 _3346_ (.A(_0409_),
    .ZN(_0410_));
 NAND2_X2 _3347_ (.A1(_0264_),
    .A2(_0410_),
    .ZN(_0411_));
 NOR2_X4 _3348_ (.A1(_0121_),
    .A2(net132),
    .ZN(_0412_));
 INV_X2 _3349_ (.A(_0412_),
    .ZN(_0413_));
 NAND3_X2 _3350_ (.A1(_0261_),
    .A2(_0263_),
    .A3(_0413_),
    .ZN(_0414_));
 NAND2_X2 _3351_ (.A1(_0411_),
    .A2(_0414_),
    .ZN(_0415_));
 NAND2_X2 _3352_ (.A1(_0415_),
    .A2(_0284_),
    .ZN(_0416_));
 NAND2_X2 _3353_ (.A1(_0408_),
    .A2(_0416_),
    .ZN(_0417_));
 INV_X2 _3354_ (.A(_0417_),
    .ZN(_0418_));
 TAPCELL_X1 PHY_40 ();
 NAND2_X1 _3356_ (.A1(_0418_),
    .A2(net104),
    .ZN(_0420_));
 TAPCELL_X1 PHY_39 ();
 NAND3_X1 _3358_ (.A1(_0400_),
    .A2(_0420_),
    .A3(net87),
    .ZN(_0422_));
 AOI21_X1 _3359_ (.A(_0344_),
    .B1(_0382_),
    .B2(_0422_),
    .ZN(_0423_));
 NOR2_X1 _3360_ (.A1(_0343_),
    .A2(_0423_),
    .ZN(_2187_));
 INV_X4 _3361_ (.A(net81),
    .ZN(_0424_));
 TAPCELL_X1 PHY_38 ();
 TAPCELL_X1 PHY_37 ();
 NAND2_X1 _3364_ (.A1(_0256_),
    .A2(_0270_),
    .ZN(_0427_));
 TAPCELL_X1 PHY_36 ();
 NAND2_X1 _3366_ (.A1(_0427_),
    .A2(_0284_),
    .ZN(_0429_));
 NAND2_X1 _3367_ (.A1(_0290_),
    .A2(_0293_),
    .ZN(_0430_));
 NAND2_X1 _3368_ (.A1(_0430_),
    .A2(_0274_),
    .ZN(_0431_));
 TAPCELL_X1 PHY_35 ();
 NAND3_X1 _3370_ (.A1(_0429_),
    .A2(_0431_),
    .A3(_0295_),
    .ZN(_0433_));
 NAND3_X1 _3371_ (.A1(_0347_),
    .A2(_0350_),
    .A3(_0284_),
    .ZN(_0434_));
 INV_X1 _3372_ (.A(_0282_),
    .ZN(_0435_));
 NAND2_X1 _3373_ (.A1(_0264_),
    .A2(_0435_),
    .ZN(_0436_));
 NAND3_X1 _3374_ (.A1(_0261_),
    .A2(_0263_),
    .A3(_0279_),
    .ZN(_0437_));
 NAND3_X1 _3375_ (.A1(_0436_),
    .A2(_0437_),
    .A3(_0274_),
    .ZN(_0438_));
 NAND3_X1 _3376_ (.A1(_0434_),
    .A2(_0438_),
    .A3(net104),
    .ZN(_0439_));
 NAND3_X1 _3377_ (.A1(_0433_),
    .A2(_0439_),
    .A3(net115),
    .ZN(_0440_));
 NAND3_X1 _3378_ (.A1(_0284_),
    .A2(_0251_),
    .A3(_0298_),
    .ZN(_0441_));
 NOR2_X1 _3379_ (.A1(_0441_),
    .A2(_0295_),
    .ZN(_0442_));
 NAND2_X1 _3380_ (.A1(_0442_),
    .A2(_0305_),
    .ZN(_0443_));
 NAND2_X1 _3381_ (.A1(_0440_),
    .A2(_0443_),
    .ZN(_0444_));
 AOI21_X1 _3382_ (.A(_0424_),
    .B1(_0444_),
    .B2(_0344_),
    .ZN(_0445_));
 INV_X1 _3383_ (.A(_0445_),
    .ZN(_0446_));
 INV_X2 _3384_ (.A(_0317_),
    .ZN(_0447_));
 NAND2_X1 _3385_ (.A1(_0397_),
    .A2(_0274_),
    .ZN(_0448_));
 NAND2_X1 _3386_ (.A1(_0407_),
    .A2(_0284_),
    .ZN(_0449_));
 NAND2_X1 _3387_ (.A1(_0448_),
    .A2(_0449_),
    .ZN(_0450_));
 NAND2_X1 _3388_ (.A1(_0450_),
    .A2(_0295_),
    .ZN(_0451_));
 TAPCELL_X1 PHY_34 ();
 NAND3_X1 _3390_ (.A1(_0325_),
    .A2(_0328_),
    .A3(_0284_),
    .ZN(_0453_));
 NAND3_X1 _3391_ (.A1(_0411_),
    .A2(_0414_),
    .A3(_0274_),
    .ZN(_0454_));
 NAND3_X1 _3392_ (.A1(_0453_),
    .A2(_0454_),
    .A3(net104),
    .ZN(_0455_));
 NAND3_X1 _3393_ (.A1(_0451_),
    .A2(net86),
    .A3(_0455_),
    .ZN(_0456_));
 NAND3_X1 _3394_ (.A1(_0363_),
    .A2(_0367_),
    .A3(_0284_),
    .ZN(_0457_));
 INV_X1 _3395_ (.A(_0356_),
    .ZN(_0458_));
 NAND2_X1 _3396_ (.A1(_0264_),
    .A2(_0458_),
    .ZN(_0459_));
 INV_X1 _3397_ (.A(_0354_),
    .ZN(_0460_));
 NAND3_X1 _3398_ (.A1(_0261_),
    .A2(_0263_),
    .A3(_0460_),
    .ZN(_0461_));
 NAND3_X1 _3399_ (.A1(_0459_),
    .A2(_0461_),
    .A3(_0274_),
    .ZN(_0462_));
 NAND3_X1 _3400_ (.A1(_0457_),
    .A2(_0462_),
    .A3(_0295_),
    .ZN(_0463_));
 NAND3_X1 _3401_ (.A1(_0385_),
    .A2(_0388_),
    .A3(_0284_),
    .ZN(_0464_));
 NAND3_X1 _3402_ (.A1(_0372_),
    .A2(_0375_),
    .A3(_0274_),
    .ZN(_0465_));
 NAND3_X1 _3403_ (.A1(_0464_),
    .A2(_0465_),
    .A3(net104),
    .ZN(_0466_));
 NAND3_X1 _3404_ (.A1(_0463_),
    .A2(_0466_),
    .A3(_0305_),
    .ZN(_0467_));
 TAPCELL_X1 PHY_33 ();
 NAND3_X1 _3406_ (.A1(_0456_),
    .A2(_0467_),
    .A3(net84),
    .ZN(_0469_));
 NAND2_X1 _3407_ (.A1(_0319_),
    .A2(_0321_),
    .ZN(_0470_));
 NAND2_X1 _3408_ (.A1(_0470_),
    .A2(_0274_),
    .ZN(_0471_));
 OAI21_X1 _3409_ (.A(_0284_),
    .B1(_0251_),
    .B2(_0332_),
    .ZN(_0472_));
 NAND3_X1 _3410_ (.A1(_0471_),
    .A2(_0295_),
    .A3(_0472_),
    .ZN(_0473_));
 TAPCELL_X1 PHY_32 ();
 OAI21_X1 _3412_ (.A(_0341_),
    .B1(_0473_),
    .B2(net87),
    .ZN(_0475_));
 NAND4_X1 _3413_ (.A1(_0446_),
    .A2(_0447_),
    .A3(_0469_),
    .A4(_0475_),
    .ZN(_0476_));
 INV_X1 _3414_ (.A(_0476_),
    .ZN(_2183_));
 TAPCELL_X1 PHY_31 ();
 NAND2_X1 _3416_ (.A1(_0360_),
    .A2(_0232_),
    .ZN(_0478_));
 TAPCELL_X1 PHY_30 ();
 NAND3_X1 _3418_ (.A1(_0276_),
    .A2(_0286_),
    .A3(_0295_),
    .ZN(_0480_));
 NAND3_X1 _3419_ (.A1(_0478_),
    .A2(net87),
    .A3(_0480_),
    .ZN(_0481_));
 NAND3_X1 _3420_ (.A1(_0294_),
    .A2(_0232_),
    .A3(_0300_),
    .ZN(_0482_));
 INV_X1 _3421_ (.A(_0482_),
    .ZN(_0483_));
 OAI21_X1 _3422_ (.A(_0481_),
    .B1(net87),
    .B2(_0483_),
    .ZN(_0484_));
 OAI21_X1 _3423_ (.A(net81),
    .B1(_0484_),
    .B2(_2120_),
    .ZN(_0485_));
 NAND2_X1 _3424_ (.A1(_0323_),
    .A2(_0330_),
    .ZN(_0486_));
 NAND3_X1 _3425_ (.A1(_0486_),
    .A2(_0230_),
    .A3(_0231_),
    .ZN(_0487_));
 TAPCELL_X1 PHY_29 ();
 NAND2_X1 _3427_ (.A1(_0418_),
    .A2(_0295_),
    .ZN(_0488_));
 NAND3_X1 _3428_ (.A1(_0487_),
    .A2(net87),
    .A3(_0488_),
    .ZN(_0489_));
 NAND2_X2 _3429_ (.A1(_0398_),
    .A2(_0232_),
    .ZN(_0490_));
 NAND3_X1 _3430_ (.A1(_0369_),
    .A2(_0377_),
    .A3(_0295_),
    .ZN(_0491_));
 NAND3_X1 _3431_ (.A1(_0490_),
    .A2(_0305_),
    .A3(_0491_),
    .ZN(_0492_));
 NAND2_X1 _3432_ (.A1(_0489_),
    .A2(_0492_),
    .ZN(_0493_));
 NAND2_X1 _3433_ (.A1(_0493_),
    .A2(_2120_),
    .ZN(_0494_));
 TAPCELL_X1 PHY_28 ();
 NOR2_X1 _3435_ (.A1(_0334_),
    .A2(net104),
    .ZN(_0496_));
 INV_X1 _3436_ (.A(_0496_),
    .ZN(_0497_));
 NOR2_X1 _3437_ (.A1(_0497_),
    .A2(net87),
    .ZN(_0498_));
 INV_X1 _3438_ (.A(_0498_),
    .ZN(_0499_));
 AOI21_X1 _3439_ (.A(_0317_),
    .B1(_0499_),
    .B2(_0341_),
    .ZN(_0500_));
 AND3_X1 _3440_ (.A1(_0485_),
    .A2(_0494_),
    .A3(_0500_),
    .ZN(_2179_));
 NAND3_X1 _3441_ (.A1(_0429_),
    .A2(_0431_),
    .A3(net104),
    .ZN(_0501_));
 NAND2_X1 _3442_ (.A1(_0441_),
    .A2(_0295_),
    .ZN(_0502_));
 NAND2_X1 _3443_ (.A1(_0501_),
    .A2(_0502_),
    .ZN(_0503_));
 NAND2_X1 _3444_ (.A1(_0503_),
    .A2(_0305_),
    .ZN(_0504_));
 TAPCELL_X1 PHY_27 ();
 NAND2_X1 _3446_ (.A1(_0368_),
    .A2(_0284_),
    .ZN(_0506_));
 NAND3_X1 _3447_ (.A1(_0355_),
    .A2(_0357_),
    .A3(_0274_),
    .ZN(_0507_));
 NAND3_X1 _3448_ (.A1(_0506_),
    .A2(_0507_),
    .A3(net104),
    .ZN(_0508_));
 NAND2_X1 _3449_ (.A1(_0351_),
    .A2(_0284_),
    .ZN(_0509_));
 NAND3_X1 _3450_ (.A1(_0281_),
    .A2(_0283_),
    .A3(_0274_),
    .ZN(_0510_));
 NAND3_X1 _3451_ (.A1(_0509_),
    .A2(_0510_),
    .A3(_0295_),
    .ZN(_0511_));
 NAND3_X1 _3452_ (.A1(_0508_),
    .A2(_0511_),
    .A3(net86),
    .ZN(_0512_));
 NAND3_X1 _3453_ (.A1(_0504_),
    .A2(_0512_),
    .A3(net81),
    .ZN(_0513_));
 NAND3_X1 _3454_ (.A1(_0448_),
    .A2(_0449_),
    .A3(net104),
    .ZN(_0514_));
 NAND2_X1 _3455_ (.A1(_0464_),
    .A2(_0465_),
    .ZN(_0515_));
 NAND2_X1 _3456_ (.A1(_0515_),
    .A2(_0295_),
    .ZN(_0516_));
 NAND3_X1 _3457_ (.A1(_0514_),
    .A2(_0516_),
    .A3(_0305_),
    .ZN(_0517_));
 NAND2_X1 _3458_ (.A1(_0325_),
    .A2(_0328_),
    .ZN(_0518_));
 NAND2_X1 _3459_ (.A1(_0518_),
    .A2(_0284_),
    .ZN(_0519_));
 NAND2_X1 _3460_ (.A1(_0415_),
    .A2(_0274_),
    .ZN(_0520_));
 NAND3_X1 _3461_ (.A1(_0519_),
    .A2(_0520_),
    .A3(_0295_),
    .ZN(_0521_));
 NAND3_X1 _3462_ (.A1(_0471_),
    .A2(net117),
    .A3(_0472_),
    .ZN(_0522_));
 NAND3_X1 _3463_ (.A1(_0521_),
    .A2(_0522_),
    .A3(net115),
    .ZN(_0523_));
 NAND3_X1 _3464_ (.A1(_0517_),
    .A2(_0523_),
    .A3(net83),
    .ZN(_0524_));
 NAND2_X1 _3465_ (.A1(_0513_),
    .A2(_0524_),
    .ZN(_0525_));
 NOR2_X1 _3466_ (.A1(_0424_),
    .A2(_0344_),
    .ZN(_0526_));
 INV_X1 _3467_ (.A(_0526_),
    .ZN(_0527_));
 NAND2_X1 _3468_ (.A1(_0527_),
    .A2(_0447_),
    .ZN(_0528_));
 INV_X1 _3469_ (.A(_0528_),
    .ZN(_0529_));
 NAND2_X1 _3470_ (.A1(_0525_),
    .A2(_0529_),
    .ZN(_0530_));
 INV_X1 _3471_ (.A(_0530_),
    .ZN(_2176_));
 NAND2_X1 _3472_ (.A1(_0302_),
    .A2(_0305_),
    .ZN(_0531_));
 OAI21_X1 _3473_ (.A(_0531_),
    .B1(_0380_),
    .B2(_0305_),
    .ZN(_0532_));
 NAND2_X1 _3474_ (.A1(_0532_),
    .A2(net81),
    .ZN(_0533_));
 NAND3_X1 _3475_ (.A1(_0400_),
    .A2(_0420_),
    .A3(_0305_),
    .ZN(_0534_));
 OAI21_X1 _3476_ (.A(_0534_),
    .B1(_0305_),
    .B2(_0337_),
    .ZN(_0535_));
 OAI21_X1 _3477_ (.A(_0533_),
    .B1(_0344_),
    .B2(_0535_),
    .ZN(_0536_));
 NAND2_X1 _3478_ (.A1(_0536_),
    .A2(_0529_),
    .ZN(_0537_));
 INV_X1 _3479_ (.A(_0537_),
    .ZN(_2172_));
 AOI21_X1 _3480_ (.A(net115),
    .B1(_0433_),
    .B2(_0439_),
    .ZN(_0538_));
 AOI21_X1 _3481_ (.A(_0305_),
    .B1(_0463_),
    .B2(_0466_),
    .ZN(_0539_));
 OR3_X1 _3482_ (.A1(_0538_),
    .A2(_0539_),
    .A3(net84),
    .ZN(_0540_));
 NAND3_X1 _3483_ (.A1(_0442_),
    .A2(net84),
    .A3(net115),
    .ZN(_0541_));
 NAND3_X1 _3484_ (.A1(_0540_),
    .A2(net81),
    .A3(_0541_),
    .ZN(_0542_));
 AOI21_X1 _3485_ (.A(_0344_),
    .B1(_0473_),
    .B2(net115),
    .ZN(_0543_));
 AND2_X1 _3486_ (.A1(_0451_),
    .A2(_0455_),
    .ZN(_0544_));
 OAI21_X1 _3487_ (.A(_0543_),
    .B1(_0544_),
    .B2(net115),
    .ZN(_0545_));
 AOI21_X1 _3488_ (.A(_0317_),
    .B1(_0545_),
    .B2(_0424_),
    .ZN(_0546_));
 NAND2_X1 _3489_ (.A1(_0542_),
    .A2(_0546_),
    .ZN(_0547_));
 INV_X1 _3490_ (.A(_0547_),
    .ZN(_2167_));
 NAND3_X1 _3491_ (.A1(_0490_),
    .A2(_0491_),
    .A3(net87),
    .ZN(_0548_));
 NAND3_X1 _3492_ (.A1(_0478_),
    .A2(_0305_),
    .A3(_0480_),
    .ZN(_0549_));
 NAND3_X1 _3493_ (.A1(_0548_),
    .A2(_0549_),
    .A3(_0344_),
    .ZN(_0550_));
 NAND3_X1 _3494_ (.A1(_0483_),
    .A2(net83),
    .A3(net87),
    .ZN(_0551_));
 NAND3_X1 _3495_ (.A1(_0550_),
    .A2(net81),
    .A3(_0551_),
    .ZN(_0552_));
 NAND3_X1 _3496_ (.A1(_0487_),
    .A2(_0305_),
    .A3(_0488_),
    .ZN(_0553_));
 AOI21_X1 _3497_ (.A(_0344_),
    .B1(_0497_),
    .B2(net87),
    .ZN(_0554_));
 NAND2_X1 _3498_ (.A1(_0553_),
    .A2(_0554_),
    .ZN(_0555_));
 AOI21_X1 _3499_ (.A(_0317_),
    .B1(_0555_),
    .B2(_0424_),
    .ZN(_0556_));
 NAND2_X1 _3500_ (.A1(_0552_),
    .A2(_0556_),
    .ZN(_0557_));
 INV_X1 _3501_ (.A(_0557_),
    .ZN(_2164_));
 NAND4_X1 _3502_ (.A1(_0501_),
    .A2(net115),
    .A3(net81),
    .A4(_0502_),
    .ZN(_0558_));
 NAND2_X1 _3503_ (.A1(_0521_),
    .A2(_0522_),
    .ZN(_0559_));
 NAND3_X1 _3504_ (.A1(_0559_),
    .A2(_0305_),
    .A3(_0424_),
    .ZN(_0560_));
 NAND2_X1 _3505_ (.A1(_0558_),
    .A2(_0560_),
    .ZN(_0561_));
 NAND2_X1 _3506_ (.A1(_0561_),
    .A2(net84),
    .ZN(_0562_));
 NAND3_X1 _3507_ (.A1(_0508_),
    .A2(_0511_),
    .A3(_0305_),
    .ZN(_0563_));
 NAND3_X1 _3508_ (.A1(_0514_),
    .A2(_0516_),
    .A3(net86),
    .ZN(_0564_));
 NOR2_X2 _3509_ (.A1(_0424_),
    .A2(net82),
    .ZN(_0565_));
 NAND3_X1 _3510_ (.A1(_0563_),
    .A2(_0564_),
    .A3(_0565_),
    .ZN(_0566_));
 NAND2_X1 _3511_ (.A1(_0562_),
    .A2(_0566_),
    .ZN(_0567_));
 NAND2_X1 _3512_ (.A1(_0567_),
    .A2(_0447_),
    .ZN(_0568_));
 INV_X1 _3513_ (.A(_0568_),
    .ZN(_2159_));
 NAND3_X1 _3514_ (.A1(_0302_),
    .A2(net87),
    .A3(net81),
    .ZN(_0569_));
 NAND4_X1 _3515_ (.A1(_0331_),
    .A2(_0305_),
    .A3(_0424_),
    .A4(_0336_),
    .ZN(_0570_));
 NAND2_X1 _3516_ (.A1(_0569_),
    .A2(_0570_),
    .ZN(_0571_));
 NAND2_X1 _3517_ (.A1(_0571_),
    .A2(_2120_),
    .ZN(_0572_));
 NAND3_X1 _3518_ (.A1(_0382_),
    .A2(_0422_),
    .A3(_0565_),
    .ZN(_0573_));
 NAND2_X1 _3519_ (.A1(_0572_),
    .A2(_0573_),
    .ZN(_0574_));
 NAND2_X1 _3520_ (.A1(_0574_),
    .A2(_0447_),
    .ZN(_0575_));
 INV_X1 _3521_ (.A(_0575_),
    .ZN(_2156_));
 NAND3_X1 _3522_ (.A1(_0456_),
    .A2(_0467_),
    .A3(_0344_),
    .ZN(_0576_));
 NAND3_X1 _3523_ (.A1(_0440_),
    .A2(net84),
    .A3(_0443_),
    .ZN(_0577_));
 NAND2_X1 _3524_ (.A1(_0576_),
    .A2(_0577_),
    .ZN(_0578_));
 NAND2_X1 _3525_ (.A1(_0578_),
    .A2(net81),
    .ZN(_0579_));
 NOR2_X1 _3526_ (.A1(_0473_),
    .A2(net87),
    .ZN(_0580_));
 NAND2_X1 _3527_ (.A1(_0580_),
    .A2(net83),
    .ZN(_0581_));
 AOI21_X1 _3528_ (.A(_0317_),
    .B1(_0581_),
    .B2(_0424_),
    .ZN(_0582_));
 AND2_X1 _3529_ (.A1(_0579_),
    .A2(_0582_),
    .ZN(_2152_));
 NAND2_X1 _3530_ (.A1(_0251_),
    .A2(_0332_),
    .ZN(_0583_));
 NAND2_X1 _3531_ (.A1(_0264_),
    .A2(_0318_),
    .ZN(_0584_));
 NAND2_X1 _3532_ (.A1(_0583_),
    .A2(_0584_),
    .ZN(_0585_));
 NOR2_X1 _3533_ (.A1(_0585_),
    .A2(_0284_),
    .ZN(_0586_));
 NAND3_X1 _3534_ (.A1(_0586_),
    .A2(_0305_),
    .A3(_0295_),
    .ZN(_0587_));
 TAPCELL_X1 PHY_26 ();
 OAI21_X1 _3536_ (.A(_0424_),
    .B1(_0587_),
    .B2(_0344_),
    .ZN(_0589_));
 NAND2_X1 _3537_ (.A1(_0589_),
    .A2(_0447_),
    .ZN(_0590_));
 NAND2_X1 _3538_ (.A1(_0251_),
    .A2(_0320_),
    .ZN(_0591_));
 NAND2_X1 _3539_ (.A1(_0264_),
    .A2(_0324_),
    .ZN(_0592_));
 NAND3_X1 _3540_ (.A1(_0591_),
    .A2(_0592_),
    .A3(_0284_),
    .ZN(_0593_));
 NAND2_X1 _3541_ (.A1(_0264_),
    .A2(_0413_),
    .ZN(_0594_));
 NAND3_X1 _3542_ (.A1(_0261_),
    .A2(_0263_),
    .A3(_0327_),
    .ZN(_0595_));
 NAND3_X1 _3543_ (.A1(_0594_),
    .A2(_0595_),
    .A3(_0274_),
    .ZN(_0596_));
 AND2_X1 _3544_ (.A1(_0593_),
    .A2(_0596_),
    .ZN(_0597_));
 INV_X1 _3545_ (.A(_0597_),
    .ZN(_0598_));
 NAND2_X1 _3546_ (.A1(_0598_),
    .A2(net114),
    .ZN(_0599_));
 NAND2_X1 _3547_ (.A1(_0251_),
    .A2(_0404_),
    .ZN(_0600_));
 NAND2_X1 _3548_ (.A1(_0264_),
    .A2(_0391_),
    .ZN(_0601_));
 NAND2_X1 _3549_ (.A1(_0600_),
    .A2(_0601_),
    .ZN(_0602_));
 INV_X1 _3550_ (.A(_0602_),
    .ZN(_0603_));
 TAPCELL_X1 PHY_25 ();
 NAND2_X1 _3552_ (.A1(_0603_),
    .A2(_0274_),
    .ZN(_0605_));
 NAND2_X1 _3553_ (.A1(_0251_),
    .A2(_0410_),
    .ZN(_0606_));
 NAND2_X1 _3554_ (.A1(_0264_),
    .A2(_0402_),
    .ZN(_0607_));
 NAND2_X1 _3555_ (.A1(_0606_),
    .A2(_0607_),
    .ZN(_0608_));
 NAND2_X1 _3556_ (.A1(_0608_),
    .A2(_0284_),
    .ZN(_0609_));
 NAND3_X1 _3557_ (.A1(_0605_),
    .A2(_0295_),
    .A3(_0609_),
    .ZN(_0610_));
 NAND3_X1 _3558_ (.A1(_0599_),
    .A2(_0610_),
    .A3(net85),
    .ZN(_0611_));
 NAND2_X1 _3559_ (.A1(_0251_),
    .A2(_0383_),
    .ZN(_0612_));
 NAND2_X1 _3560_ (.A1(_0264_),
    .A2(_0373_),
    .ZN(_0613_));
 NAND2_X1 _3561_ (.A1(_0612_),
    .A2(_0613_),
    .ZN(_0614_));
 INV_X1 _3562_ (.A(_0614_),
    .ZN(_0615_));
 NAND2_X1 _3563_ (.A1(_0615_),
    .A2(_0274_),
    .ZN(_0616_));
 NAND2_X1 _3564_ (.A1(_0251_),
    .A2(_0394_),
    .ZN(_0617_));
 NAND2_X1 _3565_ (.A1(_0264_),
    .A2(_0386_),
    .ZN(_0618_));
 NAND3_X1 _3566_ (.A1(_0617_),
    .A2(_0618_),
    .A3(_0284_),
    .ZN(_0619_));
 NAND3_X1 _3567_ (.A1(_0616_),
    .A2(_0619_),
    .A3(net114),
    .ZN(_0620_));
 NAND2_X1 _3568_ (.A1(_0251_),
    .A2(_0365_),
    .ZN(_0621_));
 NAND2_X1 _3569_ (.A1(_0264_),
    .A2(_0354_),
    .ZN(_0622_));
 NAND3_X1 _3570_ (.A1(_0621_),
    .A2(_0622_),
    .A3(_0274_),
    .ZN(_0623_));
 NAND2_X1 _3571_ (.A1(_0251_),
    .A2(_0370_),
    .ZN(_0624_));
 INV_X1 _3572_ (.A(_0362_),
    .ZN(_0625_));
 NAND2_X1 _3573_ (.A1(_0264_),
    .A2(_0625_),
    .ZN(_0626_));
 NAND3_X1 _3574_ (.A1(_0624_),
    .A2(_0626_),
    .A3(_0284_),
    .ZN(_0627_));
 NAND3_X1 _3575_ (.A1(_0623_),
    .A2(_0627_),
    .A3(_0295_),
    .ZN(_0628_));
 NAND3_X1 _3576_ (.A1(_0620_),
    .A2(_0628_),
    .A3(_0305_),
    .ZN(_0629_));
 NAND2_X1 _3577_ (.A1(_0611_),
    .A2(_0629_),
    .ZN(_0630_));
 NAND2_X1 _3578_ (.A1(_0630_),
    .A2(_0344_),
    .ZN(_0631_));
 NAND2_X1 _3579_ (.A1(_0251_),
    .A2(_0292_),
    .ZN(_0632_));
 NAND2_X1 _3580_ (.A1(_0264_),
    .A2(_0298_),
    .ZN(_0633_));
 NAND2_X1 _3581_ (.A1(_0632_),
    .A2(_0633_),
    .ZN(_0634_));
 NAND2_X1 _3582_ (.A1(_0634_),
    .A2(_0284_),
    .ZN(_0635_));
 NOR2_X1 _3583_ (.A1(_0635_),
    .A2(_0295_),
    .ZN(_0636_));
 NAND2_X1 _3584_ (.A1(_0636_),
    .A2(_0305_),
    .ZN(_0637_));
 NAND3_X1 _3585_ (.A1(_0264_),
    .A2(net99),
    .A3(_0158_),
    .ZN(_0638_));
 NAND2_X1 _3586_ (.A1(_0251_),
    .A2(_0356_),
    .ZN(_0639_));
 NAND3_X1 _3587_ (.A1(_0638_),
    .A2(_0284_),
    .A3(_0639_),
    .ZN(_0640_));
 NAND2_X1 _3588_ (.A1(_0251_),
    .A2(_0348_),
    .ZN(_0641_));
 NAND2_X1 _3589_ (.A1(_0264_),
    .A2(_0280_),
    .ZN(_0642_));
 NAND2_X1 _3590_ (.A1(_0641_),
    .A2(_0642_),
    .ZN(_0643_));
 INV_X1 _3591_ (.A(_0643_),
    .ZN(_0644_));
 NAND2_X1 _3592_ (.A1(_0644_),
    .A2(_0274_),
    .ZN(_0645_));
 NAND3_X1 _3593_ (.A1(_0640_),
    .A2(_0645_),
    .A3(_0232_),
    .ZN(_0646_));
 NAND2_X1 _3594_ (.A1(_0251_),
    .A2(_0435_),
    .ZN(_0647_));
 NAND2_X1 _3595_ (.A1(_0264_),
    .A2(_0254_),
    .ZN(_0648_));
 NAND3_X1 _3596_ (.A1(_0647_),
    .A2(_0648_),
    .A3(_0284_),
    .ZN(_0649_));
 NAND2_X1 _3597_ (.A1(_0264_),
    .A2(_0288_),
    .ZN(_0650_));
 INV_X1 _3598_ (.A(_0269_),
    .ZN(_0651_));
 NAND3_X1 _3599_ (.A1(_0261_),
    .A2(_0263_),
    .A3(_0651_),
    .ZN(_0652_));
 NAND3_X1 _3600_ (.A1(_0650_),
    .A2(_0652_),
    .A3(_0274_),
    .ZN(_0653_));
 NAND2_X1 _3601_ (.A1(_0649_),
    .A2(_0653_),
    .ZN(_0654_));
 NAND2_X1 _3602_ (.A1(_0654_),
    .A2(_0295_),
    .ZN(_0655_));
 AND2_X1 _3603_ (.A1(_0646_),
    .A2(_0655_),
    .ZN(_0656_));
 OAI21_X1 _3604_ (.A(_0637_),
    .B1(_0656_),
    .B2(_0305_),
    .ZN(_0657_));
 OAI21_X1 _3605_ (.A(_0631_),
    .B1(_0657_),
    .B2(_0344_),
    .ZN(_0658_));
 AOI21_X1 _3606_ (.A(_0590_),
    .B1(_0658_),
    .B2(net81),
    .ZN(_2149_));
 XOR2_X1 _3607_ (.A(_2053_),
    .B(_2136_),
    .Z(net67));
 NAND2_X2 _3608_ (.A1(_2134_),
    .A2(_2049_),
    .ZN(_0659_));
 INV_X1 _3609_ (.A(_2133_),
    .ZN(_0660_));
 NAND2_X2 _3610_ (.A1(_0659_),
    .A2(_0660_),
    .ZN(_0661_));
 AOI21_X4 _3611_ (.A(_2135_),
    .B1(_0661_),
    .B2(_2136_),
    .ZN(_2056_));
 XNOR2_X1 _3612_ (.A(_2058_),
    .B(_2141_),
    .ZN(net69));
 XNOR2_X1 _3613_ (.A(_2144_),
    .B(_2062_),
    .ZN(net72));
 NOR2_X2 _3614_ (.A1(_2128_),
    .A2(_2131_),
    .ZN(_0662_));
 NAND2_X4 _3615_ (.A1(_0315_),
    .A2(_0662_),
    .ZN(_0663_));
 OR2_X1 _3616_ (.A1(_0663_),
    .A2(_0095_),
    .ZN(_0664_));
 TAPCELL_X1 PHY_24 ();
 NAND2_X1 _3618_ (.A1(_0664_),
    .A2(_0251_),
    .ZN(_0666_));
 TAPCELL_X1 PHY_23 ();
 TAPCELL_X1 PHY_22 ();
 OAI21_X1 _3621_ (.A(_0264_),
    .B1(_0663_),
    .B2(_2005_),
    .ZN(_0669_));
 NAND3_X1 _3622_ (.A1(_0666_),
    .A2(_0284_),
    .A3(_0669_),
    .ZN(_0670_));
 TAPCELL_X1 PHY_21 ();
 OAI21_X1 _3624_ (.A(_0264_),
    .B1(_0663_),
    .B2(_2000_),
    .ZN(_0672_));
 NAND3_X1 _3625_ (.A1(_0315_),
    .A2(_0088_),
    .A3(_0662_),
    .ZN(_0673_));
 NAND2_X1 _3626_ (.A1(_0673_),
    .A2(_0251_),
    .ZN(_0674_));
 NAND3_X1 _3627_ (.A1(_0672_),
    .A2(_0274_),
    .A3(_0674_),
    .ZN(_0675_));
 NAND2_X1 _3628_ (.A1(_0670_),
    .A2(_0675_),
    .ZN(_0676_));
 OAI21_X1 _3629_ (.A(_0251_),
    .B1(_0663_),
    .B2(_1995_),
    .ZN(_0677_));
 OAI21_X1 _3630_ (.A(_0264_),
    .B1(_0663_),
    .B2(_0159_),
    .ZN(_0678_));
 NAND3_X1 _3631_ (.A1(_0677_),
    .A2(_0678_),
    .A3(_0274_),
    .ZN(_0679_));
 OAI21_X1 _3632_ (.A(_0251_),
    .B1(_0663_),
    .B2(_2000_),
    .ZN(_0680_));
 INV_X1 _3633_ (.A(_0160_),
    .ZN(_0681_));
 NAND3_X1 _3634_ (.A1(_0315_),
    .A2(_0681_),
    .A3(_0662_),
    .ZN(_0682_));
 NAND2_X1 _3635_ (.A1(_0682_),
    .A2(_0264_),
    .ZN(_0683_));
 NAND3_X1 _3636_ (.A1(_0680_),
    .A2(_0284_),
    .A3(_0683_),
    .ZN(_0684_));
 NAND2_X1 _3637_ (.A1(_0679_),
    .A2(_0684_),
    .ZN(_0685_));
 NOR2_X1 _3638_ (.A1(_0676_),
    .A2(_0685_),
    .ZN(_0686_));
 NAND3_X1 _3639_ (.A1(_0672_),
    .A2(_0284_),
    .A3(_0674_),
    .ZN(_0687_));
 OAI21_X1 _3640_ (.A(_0264_),
    .B1(_0663_),
    .B2(_1995_),
    .ZN(_0688_));
 NAND2_X1 _3641_ (.A1(_0682_),
    .A2(_0251_),
    .ZN(_0689_));
 NAND3_X1 _3642_ (.A1(_0688_),
    .A2(_0274_),
    .A3(_0689_),
    .ZN(_0690_));
 NAND2_X1 _3643_ (.A1(_0687_),
    .A2(_0690_),
    .ZN(_0691_));
 OAI21_X1 _3644_ (.A(_0251_),
    .B1(_0663_),
    .B2(_2005_),
    .ZN(_0692_));
 NAND2_X1 _3645_ (.A1(_0673_),
    .A2(_0264_),
    .ZN(_0693_));
 NAND3_X1 _3646_ (.A1(_0692_),
    .A2(_0284_),
    .A3(_0693_),
    .ZN(_0694_));
 NAND3_X1 _3647_ (.A1(_0680_),
    .A2(_0274_),
    .A3(_0683_),
    .ZN(_0695_));
 NAND2_X1 _3648_ (.A1(_0694_),
    .A2(_0695_),
    .ZN(_0696_));
 NOR2_X1 _3649_ (.A1(_0691_),
    .A2(_0696_),
    .ZN(_0697_));
 NAND2_X1 _3650_ (.A1(_0686_),
    .A2(_0697_),
    .ZN(_0698_));
 NAND2_X1 _3651_ (.A1(_0698_),
    .A2(net104),
    .ZN(_0699_));
 NOR2_X1 _3652_ (.A1(_0663_),
    .A2(_0166_),
    .ZN(_0700_));
 NAND2_X1 _3653_ (.A1(_0700_),
    .A2(_0264_),
    .ZN(_0701_));
 INV_X2 _3654_ (.A(_0663_),
    .ZN(_0702_));
 NAND3_X1 _3655_ (.A1(_0702_),
    .A2(_0070_),
    .A3(_0251_),
    .ZN(_0703_));
 NAND2_X1 _3656_ (.A1(_0701_),
    .A2(_0703_),
    .ZN(_0704_));
 NAND4_X1 _3657_ (.A1(_0315_),
    .A2(_0079_),
    .A3(_0251_),
    .A4(_0662_),
    .ZN(_0705_));
 NAND4_X1 _3658_ (.A1(_0315_),
    .A2(_0070_),
    .A3(_0264_),
    .A4(_0662_),
    .ZN(_0706_));
 NAND2_X1 _3659_ (.A1(_0705_),
    .A2(_0706_),
    .ZN(_0707_));
 NOR2_X1 _3660_ (.A1(_0704_),
    .A2(_0707_),
    .ZN(_0708_));
 NOR2_X1 _3661_ (.A1(_0663_),
    .A2(_0082_),
    .ZN(_0709_));
 NAND2_X1 _3662_ (.A1(_0709_),
    .A2(_0251_),
    .ZN(_0710_));
 NAND3_X1 _3663_ (.A1(_0702_),
    .A2(_0080_),
    .A3(_0264_),
    .ZN(_0711_));
 NAND2_X1 _3664_ (.A1(_0710_),
    .A2(_0711_),
    .ZN(_0712_));
 TAPCELL_X1 PHY_20 ();
 NAND2_X1 _3666_ (.A1(_0712_),
    .A2(_0284_),
    .ZN(_0714_));
 TAPCELL_X1 PHY_19 ();
 OAI21_X1 _3668_ (.A(_0251_),
    .B1(_0663_),
    .B2(_1985_),
    .ZN(_0716_));
 TAPCELL_X1 PHY_18 ();
 OAI21_X1 _3670_ (.A(_0264_),
    .B1(_0663_),
    .B2(_0173_),
    .ZN(_0718_));
 NAND3_X1 _3671_ (.A1(_0716_),
    .A2(_0718_),
    .A3(_0284_),
    .ZN(_0719_));
 NAND3_X1 _3672_ (.A1(_0708_),
    .A2(_0714_),
    .A3(_0719_),
    .ZN(_0720_));
 NAND2_X1 _3673_ (.A1(_0700_),
    .A2(_0251_),
    .ZN(_0721_));
 NOR2_X1 _3674_ (.A1(_0663_),
    .A2(_1975_),
    .ZN(_0722_));
 NAND2_X1 _3675_ (.A1(_0722_),
    .A2(_0251_),
    .ZN(_0723_));
 NAND2_X1 _3676_ (.A1(_0721_),
    .A2(_0723_),
    .ZN(_0724_));
 NAND2_X1 _3677_ (.A1(_0722_),
    .A2(_0264_),
    .ZN(_0725_));
 INV_X1 _3678_ (.A(_0076_),
    .ZN(_0726_));
 NAND3_X1 _3679_ (.A1(_0702_),
    .A2(_0726_),
    .A3(_0264_),
    .ZN(_0727_));
 NAND2_X1 _3680_ (.A1(_0725_),
    .A2(_0727_),
    .ZN(_0728_));
 NOR2_X1 _3681_ (.A1(_0724_),
    .A2(_0728_),
    .ZN(_0729_));
 NOR2_X1 _3682_ (.A1(_0729_),
    .A2(_0284_),
    .ZN(_0730_));
 OAI21_X1 _3683_ (.A(_0295_),
    .B1(_0720_),
    .B2(_0730_),
    .ZN(_0731_));
 NAND3_X1 _3684_ (.A1(_0710_),
    .A2(_0711_),
    .A3(_0274_),
    .ZN(_0732_));
 NOR2_X1 _3685_ (.A1(_0663_),
    .A2(_1990_),
    .ZN(_0733_));
 NAND2_X1 _3686_ (.A1(_0733_),
    .A2(_0264_),
    .ZN(_0734_));
 NAND3_X1 _3687_ (.A1(_0702_),
    .A2(_0158_),
    .A3(_0251_),
    .ZN(_0735_));
 NAND3_X1 _3688_ (.A1(_0734_),
    .A2(_0735_),
    .A3(_0284_),
    .ZN(_0736_));
 NAND2_X1 _3689_ (.A1(_0732_),
    .A2(_0736_),
    .ZN(_0737_));
 NAND2_X1 _3690_ (.A1(_0709_),
    .A2(_0264_),
    .ZN(_0738_));
 NAND2_X1 _3691_ (.A1(_0733_),
    .A2(_0251_),
    .ZN(_0739_));
 NAND2_X1 _3692_ (.A1(_0738_),
    .A2(_0739_),
    .ZN(_0740_));
 NAND2_X1 _3693_ (.A1(_0740_),
    .A2(_0284_),
    .ZN(_0741_));
 TAPCELL_X1 PHY_17 ();
 NAND3_X1 _3695_ (.A1(_0716_),
    .A2(_0718_),
    .A3(_0274_),
    .ZN(_0743_));
 NAND3_X1 _3696_ (.A1(_0737_),
    .A2(_0741_),
    .A3(_0743_),
    .ZN(_0744_));
 NAND3_X1 _3697_ (.A1(_0734_),
    .A2(_0735_),
    .A3(_0274_),
    .ZN(_0745_));
 NAND2_X1 _3698_ (.A1(_0688_),
    .A2(_0689_),
    .ZN(_0746_));
 NAND2_X1 _3699_ (.A1(_0746_),
    .A2(_0284_),
    .ZN(_0747_));
 NAND2_X1 _3700_ (.A1(_0745_),
    .A2(_0747_),
    .ZN(_0748_));
 NAND3_X1 _3701_ (.A1(_0677_),
    .A2(_0678_),
    .A3(_0284_),
    .ZN(_0749_));
 NAND2_X1 _3702_ (.A1(_0740_),
    .A2(_0274_),
    .ZN(_0750_));
 NAND3_X1 _3703_ (.A1(_0748_),
    .A2(_0749_),
    .A3(_0750_),
    .ZN(_0751_));
 NOR2_X1 _3704_ (.A1(_0744_),
    .A2(_0751_),
    .ZN(_0752_));
 NAND3_X1 _3705_ (.A1(_0699_),
    .A2(_0731_),
    .A3(_0752_),
    .ZN(_0753_));
 NAND2_X1 _3706_ (.A1(_0753_),
    .A2(_0305_),
    .ZN(_0754_));
 OR2_X1 _3707_ (.A1(_0663_),
    .A2(_2010_),
    .ZN(_0755_));
 NAND2_X1 _3708_ (.A1(_0755_),
    .A2(_0251_),
    .ZN(_0756_));
 NAND2_X1 _3709_ (.A1(_0664_),
    .A2(_0264_),
    .ZN(_0757_));
 NAND3_X1 _3710_ (.A1(_0756_),
    .A2(_0757_),
    .A3(_0274_),
    .ZN(_0758_));
 OR2_X1 _3711_ (.A1(_0663_),
    .A2(_2015_),
    .ZN(_0759_));
 NAND2_X1 _3712_ (.A1(_0759_),
    .A2(_0251_),
    .ZN(_0760_));
 OR2_X1 _3713_ (.A1(_0663_),
    .A2(_0146_),
    .ZN(_0761_));
 NAND2_X1 _3714_ (.A1(_0761_),
    .A2(_0264_),
    .ZN(_0762_));
 NAND2_X1 _3715_ (.A1(_0760_),
    .A2(_0762_),
    .ZN(_0763_));
 OAI21_X1 _3716_ (.A(_0758_),
    .B1(_0274_),
    .B2(_0763_),
    .ZN(_0764_));
 NAND2_X1 _3717_ (.A1(_0755_),
    .A2(_0264_),
    .ZN(_0765_));
 NAND2_X1 _3718_ (.A1(_0761_),
    .A2(_0251_),
    .ZN(_0766_));
 NAND3_X1 _3719_ (.A1(_0765_),
    .A2(_0766_),
    .A3(_0284_),
    .ZN(_0767_));
 NAND3_X1 _3720_ (.A1(_0666_),
    .A2(_0274_),
    .A3(_0669_),
    .ZN(_0768_));
 NAND2_X1 _3721_ (.A1(_0767_),
    .A2(_0768_),
    .ZN(_0769_));
 NOR2_X1 _3722_ (.A1(_0764_),
    .A2(_0769_),
    .ZN(_0770_));
 NAND3_X1 _3723_ (.A1(_0765_),
    .A2(_0766_),
    .A3(_0274_),
    .ZN(_0771_));
 OR2_X1 _3724_ (.A1(_0663_),
    .A2(_0127_),
    .ZN(_0772_));
 NAND2_X1 _3725_ (.A1(_0772_),
    .A2(_0251_),
    .ZN(_0773_));
 NAND2_X1 _3726_ (.A1(_0759_),
    .A2(_0264_),
    .ZN(_0774_));
 NAND2_X1 _3727_ (.A1(_0773_),
    .A2(_0774_),
    .ZN(_0775_));
 OAI21_X1 _3728_ (.A(_0771_),
    .B1(_0274_),
    .B2(_0775_),
    .ZN(_0776_));
 NAND3_X1 _3729_ (.A1(_0756_),
    .A2(_0757_),
    .A3(_0284_),
    .ZN(_0777_));
 NAND3_X1 _3730_ (.A1(_0692_),
    .A2(_0274_),
    .A3(_0693_),
    .ZN(_0778_));
 NAND2_X1 _3731_ (.A1(_0777_),
    .A2(_0778_),
    .ZN(_0779_));
 NOR2_X1 _3732_ (.A1(_0776_),
    .A2(_0779_),
    .ZN(_0780_));
 NAND2_X1 _3733_ (.A1(_0770_),
    .A2(_0780_),
    .ZN(_0781_));
 NAND3_X1 _3734_ (.A1(_0686_),
    .A2(_0697_),
    .A3(_0295_),
    .ZN(_0782_));
 NAND3_X1 _3735_ (.A1(_0763_),
    .A2(_0775_),
    .A3(_0274_),
    .ZN(_0783_));
 OR2_X1 _3736_ (.A1(_0663_),
    .A2(_0116_),
    .ZN(_0784_));
 NAND2_X1 _3737_ (.A1(_0784_),
    .A2(_0264_),
    .ZN(_0785_));
 NAND2_X1 _3738_ (.A1(_0702_),
    .A2(_0148_),
    .ZN(_0786_));
 NAND2_X1 _3739_ (.A1(_0786_),
    .A2(_0251_),
    .ZN(_0787_));
 NAND2_X1 _3740_ (.A1(_0785_),
    .A2(_0787_),
    .ZN(_0788_));
 OR2_X1 _3741_ (.A1(_0663_),
    .A2(_0121_),
    .ZN(_0789_));
 NAND2_X1 _3742_ (.A1(_0789_),
    .A2(_0251_),
    .ZN(_0790_));
 NAND2_X1 _3743_ (.A1(_0786_),
    .A2(_0264_),
    .ZN(_0791_));
 NAND2_X1 _3744_ (.A1(_0790_),
    .A2(_0791_),
    .ZN(_0792_));
 NAND3_X1 _3745_ (.A1(_0788_),
    .A2(_0792_),
    .A3(_0284_),
    .ZN(_0793_));
 NAND2_X1 _3746_ (.A1(_0783_),
    .A2(_0793_),
    .ZN(_0794_));
 NOR2_X1 _3747_ (.A1(_0663_),
    .A2(_2020_),
    .ZN(_0795_));
 NAND2_X1 _3748_ (.A1(_0772_),
    .A2(_0264_),
    .ZN(_0796_));
 NAND2_X1 _3749_ (.A1(_0784_),
    .A2(_0251_),
    .ZN(_0797_));
 AOI21_X1 _3750_ (.A(_0795_),
    .B1(_0796_),
    .B2(_0797_),
    .ZN(_0798_));
 NAND3_X1 _3751_ (.A1(_0794_),
    .A2(net104),
    .A3(_0798_),
    .ZN(_0799_));
 AOI21_X1 _3752_ (.A(_0781_),
    .B1(_0782_),
    .B2(_0799_),
    .ZN(_0800_));
 NAND2_X1 _3753_ (.A1(_0754_),
    .A2(_0800_),
    .ZN(_0801_));
 NAND2_X1 _3754_ (.A1(_0801_),
    .A2(net84),
    .ZN(_0802_));
 NAND2_X1 _3755_ (.A1(_0702_),
    .A2(_2038_),
    .ZN(_0803_));
 OAI22_X1 _3756_ (.A1(_0803_),
    .A2(_0251_),
    .B1(_0141_),
    .B2(_0663_),
    .ZN(_0804_));
 NOR2_X1 _3757_ (.A1(_0663_),
    .A2(_0136_),
    .ZN(_0805_));
 NAND2_X1 _3758_ (.A1(_0805_),
    .A2(_0264_),
    .ZN(_0806_));
 NAND2_X1 _3759_ (.A1(_0702_),
    .A2(_2035_),
    .ZN(_0807_));
 OAI211_X2 _3760_ (.A(_0806_),
    .B(_0807_),
    .C1(_0803_),
    .C2(_0264_),
    .ZN(_0808_));
 AOI21_X1 _3761_ (.A(_0804_),
    .B1(_0808_),
    .B2(_0274_),
    .ZN(_0809_));
 NOR2_X1 _3762_ (.A1(_0809_),
    .A2(net104),
    .ZN(_0810_));
 AND2_X1 _3763_ (.A1(_0808_),
    .A2(_0284_),
    .ZN(_0811_));
 AOI21_X1 _3764_ (.A(_0284_),
    .B1(_0788_),
    .B2(_0792_),
    .ZN(_0812_));
 NAND2_X1 _3765_ (.A1(_0805_),
    .A2(_0251_),
    .ZN(_0813_));
 OAI21_X1 _3766_ (.A(_0813_),
    .B1(_2030_),
    .B2(_0663_),
    .ZN(_0814_));
 NOR2_X1 _3767_ (.A1(_0789_),
    .A2(_0251_),
    .ZN(_0815_));
 OR2_X1 _3768_ (.A1(_0814_),
    .A2(_0815_),
    .ZN(_0816_));
 NOR3_X1 _3769_ (.A1(_0811_),
    .A2(_0812_),
    .A3(_0816_),
    .ZN(_0817_));
 OR2_X1 _3770_ (.A1(_0809_),
    .A2(_0295_),
    .ZN(_0818_));
 NAND2_X1 _3771_ (.A1(_0794_),
    .A2(_0798_),
    .ZN(_0819_));
 NAND2_X1 _3772_ (.A1(_0819_),
    .A2(_0295_),
    .ZN(_0820_));
 NAND3_X1 _3773_ (.A1(_0817_),
    .A2(_0818_),
    .A3(_0820_),
    .ZN(_0821_));
 NAND2_X1 _3774_ (.A1(_0344_),
    .A2(net115),
    .ZN(_0822_));
 AOI21_X1 _3775_ (.A(_0810_),
    .B1(_0821_),
    .B2(_0822_),
    .ZN(_0823_));
 NAND2_X1 _3776_ (.A1(_0802_),
    .A2(_0823_),
    .ZN(_0824_));
 NOR2_X1 _3777_ (.A1(_0317_),
    .A2(net120),
    .ZN(_0825_));
 INV_X1 _3778_ (.A(_0825_),
    .ZN(_0826_));
 NAND3_X1 _3779_ (.A1(_0274_),
    .A2(_0264_),
    .A3(_2113_),
    .ZN(_0827_));
 NOR3_X1 _3780_ (.A1(_0527_),
    .A2(_0826_),
    .A3(_0827_),
    .ZN(_0828_));
 OR3_X1 _3781_ (.A1(_0828_),
    .A2(_0424_),
    .A3(_0826_),
    .ZN(_0829_));
 INV_X1 _3782_ (.A(_0829_),
    .ZN(_0830_));
 NAND2_X1 _3783_ (.A1(_0824_),
    .A2(_0830_),
    .ZN(_0831_));
 NOR2_X1 _3784_ (.A1(_0424_),
    .A2(_0317_),
    .ZN(_0832_));
 INV_X1 _3785_ (.A(_0832_),
    .ZN(_0833_));
 NAND3_X1 _3786_ (.A1(_0649_),
    .A2(_0653_),
    .A3(net104),
    .ZN(_0834_));
 NAND2_X1 _3787_ (.A1(_0635_),
    .A2(_0295_),
    .ZN(_0835_));
 NAND2_X1 _3788_ (.A1(_0834_),
    .A2(_0835_),
    .ZN(_0836_));
 NAND2_X1 _3789_ (.A1(_0836_),
    .A2(_0305_),
    .ZN(_0837_));
 NAND3_X1 _3790_ (.A1(_0640_),
    .A2(_0645_),
    .A3(_0295_),
    .ZN(_0838_));
 NAND3_X1 _3791_ (.A1(_0623_),
    .A2(_0627_),
    .A3(net117),
    .ZN(_0839_));
 NAND3_X1 _3792_ (.A1(_0838_),
    .A2(net86),
    .A3(_0839_),
    .ZN(_0840_));
 AOI21_X1 _3793_ (.A(_0532_),
    .B1(_0837_),
    .B2(_0840_),
    .ZN(_0841_));
 AOI21_X1 _3794_ (.A(_0344_),
    .B1(_0504_),
    .B2(_0512_),
    .ZN(_0842_));
 AOI21_X1 _3795_ (.A(_0833_),
    .B1(_0841_),
    .B2(_0842_),
    .ZN(_0843_));
 AOI21_X1 _3796_ (.A(net83),
    .B1(_0517_),
    .B2(_0523_),
    .ZN(_0844_));
 NAND3_X1 _3797_ (.A1(_0605_),
    .A2(net104),
    .A3(_0609_),
    .ZN(_0845_));
 NAND3_X1 _3798_ (.A1(_0616_),
    .A2(_0619_),
    .A3(_0295_),
    .ZN(_0846_));
 NAND3_X1 _3799_ (.A1(_0845_),
    .A2(_0846_),
    .A3(_0305_),
    .ZN(_0847_));
 NAND3_X1 _3800_ (.A1(_0593_),
    .A2(_0596_),
    .A3(_0295_),
    .ZN(_0848_));
 OAI21_X1 _3801_ (.A(net104),
    .B1(_0585_),
    .B2(_0284_),
    .ZN(_0849_));
 NAND2_X1 _3802_ (.A1(_0848_),
    .A2(_0849_),
    .ZN(_0850_));
 INV_X1 _3803_ (.A(_0850_),
    .ZN(_0851_));
 OAI21_X1 _3804_ (.A(_0847_),
    .B1(_0305_),
    .B2(_0851_),
    .ZN(_0852_));
 NAND3_X1 _3805_ (.A1(_0535_),
    .A2(_0844_),
    .A3(_0852_),
    .ZN(_0853_));
 NOR3_X1 _3806_ (.A1(_0089_),
    .A2(_0161_),
    .A3(_2035_),
    .ZN(_0854_));
 NAND4_X1 _3807_ (.A1(_0854_),
    .A2(_0146_),
    .A3(_0136_),
    .A4(_0116_),
    .ZN(_0855_));
 NOR4_X1 _3808_ (.A1(_0855_),
    .A2(_0079_),
    .A3(_0158_),
    .A4(_0088_),
    .ZN(_0856_));
 NOR4_X1 _3809_ (.A1(_0726_),
    .A2(_0171_),
    .A3(_0096_),
    .A4(_0108_),
    .ZN(_0857_));
 NAND4_X1 _3810_ (.A1(_1975_),
    .A2(_2015_),
    .A3(_2025_),
    .A4(_1985_),
    .ZN(_0858_));
 NOR3_X1 _3811_ (.A1(_0128_),
    .A2(_0858_),
    .A3(_0142_),
    .ZN(_0859_));
 NOR2_X1 _3812_ (.A1(_0083_),
    .A2(_0122_),
    .ZN(_0860_));
 NAND4_X2 _3813_ (.A1(_0856_),
    .A2(_0857_),
    .A3(_0859_),
    .A4(_0860_),
    .ZN(_0861_));
 AOI22_X1 _3814_ (.A1(_0843_),
    .A2(_0853_),
    .B1(_0828_),
    .B2(_0861_),
    .ZN(_0862_));
 NAND2_X1 _3815_ (.A1(_0831_),
    .A2(_0862_),
    .ZN(_0863_));
 MUX2_X1 _3816_ (.A(_0493_),
    .B(_0484_),
    .S(net83),
    .Z(_0864_));
 NAND2_X2 _3817_ (.A1(net81),
    .A2(_0864_),
    .ZN(_0865_));
 OAI21_X1 _3818_ (.A(_0424_),
    .B1(_0499_),
    .B2(_0344_),
    .ZN(_0866_));
 NAND3_X4 _3819_ (.A1(_0865_),
    .A2(_0447_),
    .A3(_0866_),
    .ZN(_0867_));
 NAND2_X1 _3820_ (.A1(_0603_),
    .A2(_0284_),
    .ZN(_0868_));
 NAND3_X1 _3821_ (.A1(_0617_),
    .A2(_0618_),
    .A3(_0274_),
    .ZN(_0869_));
 NAND3_X1 _3822_ (.A1(_0868_),
    .A2(net114),
    .A3(_0869_),
    .ZN(_0870_));
 NAND2_X1 _3823_ (.A1(_0615_),
    .A2(_0284_),
    .ZN(_0871_));
 NAND3_X1 _3824_ (.A1(_0624_),
    .A2(_0626_),
    .A3(_0274_),
    .ZN(_0872_));
 NAND3_X1 _3825_ (.A1(_0871_),
    .A2(_0295_),
    .A3(_0872_),
    .ZN(_0873_));
 NAND3_X1 _3826_ (.A1(_0870_),
    .A2(_0873_),
    .A3(_0305_),
    .ZN(_0874_));
 NAND2_X1 _3827_ (.A1(_0591_),
    .A2(_0592_),
    .ZN(_0875_));
 NAND2_X1 _3828_ (.A1(_0875_),
    .A2(_0274_),
    .ZN(_0876_));
 NAND2_X1 _3829_ (.A1(_0585_),
    .A2(_0284_),
    .ZN(_0877_));
 NAND2_X1 _3830_ (.A1(_0876_),
    .A2(_0877_),
    .ZN(_0878_));
 NAND2_X1 _3831_ (.A1(_0878_),
    .A2(net104),
    .ZN(_0879_));
 NAND2_X1 _3832_ (.A1(_0608_),
    .A2(_0274_),
    .ZN(_0880_));
 NAND2_X1 _3833_ (.A1(_0251_),
    .A2(_0326_),
    .ZN(_0881_));
 NAND2_X1 _3834_ (.A1(_0264_),
    .A2(_0412_),
    .ZN(_0882_));
 NAND3_X1 _3835_ (.A1(_0881_),
    .A2(_0882_),
    .A3(_0284_),
    .ZN(_0883_));
 NAND2_X1 _3836_ (.A1(_0880_),
    .A2(_0883_),
    .ZN(_0884_));
 NAND2_X1 _3837_ (.A1(_0884_),
    .A2(_0295_),
    .ZN(_0885_));
 AND2_X1 _3838_ (.A1(_0879_),
    .A2(_0885_),
    .ZN(_0886_));
 OAI21_X1 _3839_ (.A(_0874_),
    .B1(_0886_),
    .B2(_0305_),
    .ZN(_0887_));
 NAND2_X1 _3840_ (.A1(_0887_),
    .A2(_0344_),
    .ZN(_0888_));
 NAND3_X1 _3841_ (.A1(_0638_),
    .A2(_0274_),
    .A3(_0639_),
    .ZN(_0889_));
 NAND3_X1 _3842_ (.A1(_0621_),
    .A2(_0622_),
    .A3(_0284_),
    .ZN(_0890_));
 NAND3_X1 _3843_ (.A1(_0889_),
    .A2(_0232_),
    .A3(_0890_),
    .ZN(_0891_));
 NAND2_X1 _3844_ (.A1(_0644_),
    .A2(_0284_),
    .ZN(_0892_));
 NAND2_X1 _3845_ (.A1(_0647_),
    .A2(_0648_),
    .ZN(_0893_));
 NAND2_X1 _3846_ (.A1(_0893_),
    .A2(_0274_),
    .ZN(_0894_));
 NAND3_X1 _3847_ (.A1(_0892_),
    .A2(_0295_),
    .A3(_0894_),
    .ZN(_0895_));
 NAND3_X1 _3848_ (.A1(_0891_),
    .A2(_0895_),
    .A3(net85),
    .ZN(_0896_));
 NAND2_X1 _3849_ (.A1(_0634_),
    .A2(_0274_),
    .ZN(_0897_));
 NAND3_X1 _3850_ (.A1(_0650_),
    .A2(_0652_),
    .A3(_0284_),
    .ZN(_0898_));
 AOI21_X1 _3851_ (.A(_0295_),
    .B1(_0897_),
    .B2(_0898_),
    .ZN(_0899_));
 OAI21_X1 _3852_ (.A(_0896_),
    .B1(net87),
    .B2(_0899_),
    .ZN(_0900_));
 NAND2_X1 _3853_ (.A1(_0900_),
    .A2(net83),
    .ZN(_0901_));
 NAND3_X1 _3854_ (.A1(_0888_),
    .A2(_0901_),
    .A3(_0832_),
    .ZN(_0902_));
 INV_X1 _3855_ (.A(_0902_),
    .ZN(_0903_));
 NAND3_X1 _3856_ (.A1(_0863_),
    .A2(_0867_),
    .A3(_0903_),
    .ZN(_0904_));
 OR2_X1 _3857_ (.A1(_0867_),
    .A2(_0903_),
    .ZN(_0905_));
 NAND2_X1 _3858_ (.A1(_0904_),
    .A2(_0905_),
    .ZN(_0906_));
 OAI22_X1 _3859_ (.A1(_0887_),
    .A2(_0344_),
    .B1(_0900_),
    .B2(_0424_),
    .ZN(_0907_));
 NAND2_X1 _3860_ (.A1(_0907_),
    .A2(_0529_),
    .ZN(_0908_));
 NOR2_X1 _3861_ (.A1(_0908_),
    .A2(_0530_),
    .ZN(_0909_));
 NAND3_X1 _3862_ (.A1(_0840_),
    .A2(_0837_),
    .A3(net81),
    .ZN(_0910_));
 OAI21_X1 _3863_ (.A(_0910_),
    .B1(_0852_),
    .B2(_0344_),
    .ZN(_0911_));
 NAND2_X1 _3864_ (.A1(_0911_),
    .A2(_0529_),
    .ZN(_0912_));
 NOR2_X1 _3865_ (.A1(_0537_),
    .A2(_0912_),
    .ZN(_0913_));
 NAND2_X1 _3866_ (.A1(_0909_),
    .A2(_0913_),
    .ZN(_0914_));
 NAND3_X1 _3867_ (.A1(_0889_),
    .A2(_0295_),
    .A3(_0890_),
    .ZN(_0915_));
 NAND3_X1 _3868_ (.A1(_0871_),
    .A2(net114),
    .A3(_0872_),
    .ZN(_0916_));
 NAND3_X1 _3869_ (.A1(_0915_),
    .A2(_0916_),
    .A3(net85),
    .ZN(_0917_));
 NAND3_X1 _3870_ (.A1(_0892_),
    .A2(net117),
    .A3(_0894_),
    .ZN(_0918_));
 NAND2_X1 _3871_ (.A1(_0897_),
    .A2(_0898_),
    .ZN(_0919_));
 NAND2_X1 _3872_ (.A1(_0919_),
    .A2(_0295_),
    .ZN(_0920_));
 NAND3_X1 _3873_ (.A1(_0918_),
    .A2(_0920_),
    .A3(_0305_),
    .ZN(_0921_));
 NAND3_X1 _3874_ (.A1(_0917_),
    .A2(_0921_),
    .A3(net81),
    .ZN(_0922_));
 NAND3_X1 _3875_ (.A1(_0868_),
    .A2(_0295_),
    .A3(_0869_),
    .ZN(_0923_));
 NAND3_X1 _3876_ (.A1(_0880_),
    .A2(_0883_),
    .A3(net114),
    .ZN(_0924_));
 NAND3_X1 _3877_ (.A1(_0923_),
    .A2(_0924_),
    .A3(_0305_),
    .ZN(_0925_));
 OAI21_X1 _3878_ (.A(net86),
    .B1(_0878_),
    .B2(net104),
    .ZN(_0926_));
 NAND2_X1 _3879_ (.A1(_0925_),
    .A2(_0926_),
    .ZN(_0927_));
 OAI21_X1 _3880_ (.A(_0922_),
    .B1(_0344_),
    .B2(_0927_),
    .ZN(_0928_));
 NAND2_X1 _3881_ (.A1(_0928_),
    .A2(_0529_),
    .ZN(_0929_));
 OR2_X1 _3882_ (.A1(_0547_),
    .A2(_0929_),
    .ZN(_0930_));
 NAND3_X1 _3883_ (.A1(_0646_),
    .A2(_0655_),
    .A3(_0305_),
    .ZN(_0931_));
 NAND3_X1 _3884_ (.A1(_0620_),
    .A2(_0628_),
    .A3(net85),
    .ZN(_0932_));
 NAND3_X1 _3885_ (.A1(_0931_),
    .A2(_0932_),
    .A3(_0344_),
    .ZN(_0933_));
 NAND3_X1 _3886_ (.A1(_0636_),
    .A2(net82),
    .A3(net86),
    .ZN(_0934_));
 NAND3_X1 _3887_ (.A1(_0933_),
    .A2(net81),
    .A3(_0934_),
    .ZN(_0935_));
 NAND3_X1 _3888_ (.A1(_0599_),
    .A2(_0610_),
    .A3(_0305_),
    .ZN(_0936_));
 NAND2_X1 _3889_ (.A1(_0586_),
    .A2(_0295_),
    .ZN(_0937_));
 AOI21_X1 _3890_ (.A(_0344_),
    .B1(_0937_),
    .B2(net86),
    .ZN(_0938_));
 NAND2_X1 _3891_ (.A1(_0936_),
    .A2(_0938_),
    .ZN(_0939_));
 AOI21_X1 _3892_ (.A(_0317_),
    .B1(_0939_),
    .B2(_0424_),
    .ZN(_0940_));
 NAND2_X1 _3893_ (.A1(_0935_),
    .A2(_0940_),
    .ZN(_0941_));
 NOR2_X1 _3894_ (.A1(_0557_),
    .A2(_0941_),
    .ZN(_0942_));
 INV_X1 _3895_ (.A(_0942_),
    .ZN(_0943_));
 NOR3_X1 _3896_ (.A1(_0914_),
    .A2(_0930_),
    .A3(_0943_),
    .ZN(_0944_));
 NAND3_X2 _3897_ (.A1(_0579_),
    .A2(_2150_),
    .A3(_0582_),
    .ZN(_0945_));
 NAND2_X1 _3898_ (.A1(_0918_),
    .A2(_0920_),
    .ZN(_0946_));
 NAND3_X1 _3899_ (.A1(_0946_),
    .A2(net86),
    .A3(net81),
    .ZN(_0947_));
 NAND4_X1 _3900_ (.A1(_0876_),
    .A2(_0877_),
    .A3(_0305_),
    .A4(_0295_),
    .ZN(_0948_));
 OR2_X1 _3901_ (.A1(_0948_),
    .A2(net81),
    .ZN(_0949_));
 NAND2_X1 _3902_ (.A1(_0947_),
    .A2(_0949_),
    .ZN(_0950_));
 NAND2_X1 _3903_ (.A1(_0950_),
    .A2(net82),
    .ZN(_0951_));
 NAND3_X1 _3904_ (.A1(_0915_),
    .A2(_0916_),
    .A3(_0305_),
    .ZN(_0952_));
 NAND3_X1 _3905_ (.A1(_0923_),
    .A2(_0924_),
    .A3(net85),
    .ZN(_0953_));
 AND2_X1 _3906_ (.A1(_0952_),
    .A2(_0953_),
    .ZN(_0954_));
 NAND2_X1 _3907_ (.A1(_0954_),
    .A2(_0565_),
    .ZN(_0955_));
 NAND2_X1 _3908_ (.A1(_0951_),
    .A2(_0955_),
    .ZN(_0956_));
 NAND2_X1 _3909_ (.A1(_0956_),
    .A2(_0447_),
    .ZN(_0957_));
 NOR2_X4 _3910_ (.A1(_0957_),
    .A2(_0945_),
    .ZN(_2155_));
 NAND3_X1 _3911_ (.A1(_0891_),
    .A2(_0895_),
    .A3(_0305_),
    .ZN(_0958_));
 NAND3_X1 _3912_ (.A1(_0870_),
    .A2(_0873_),
    .A3(net85),
    .ZN(_0959_));
 NAND2_X1 _3913_ (.A1(_0958_),
    .A2(_0959_),
    .ZN(_0960_));
 OAI21_X1 _3914_ (.A(_0344_),
    .B1(_0960_),
    .B2(_0424_),
    .ZN(_0961_));
 AND2_X1 _3915_ (.A1(_0899_),
    .A2(net87),
    .ZN(_0962_));
 OAI21_X1 _3916_ (.A(_0447_),
    .B1(_0962_),
    .B2(_0527_),
    .ZN(_0963_));
 AOI21_X1 _3917_ (.A(net81),
    .B1(_0886_),
    .B2(_0305_),
    .ZN(_0964_));
 NOR2_X1 _3918_ (.A1(_0963_),
    .A2(_0964_),
    .ZN(_0965_));
 NAND2_X1 _3919_ (.A1(_0961_),
    .A2(_0965_),
    .ZN(_0966_));
 NOR2_X1 _3920_ (.A1(_0568_),
    .A2(_0966_),
    .ZN(_0967_));
 NAND4_X1 _3921_ (.A1(_0848_),
    .A2(_0849_),
    .A3(_0305_),
    .A4(_0424_),
    .ZN(_0968_));
 NAND4_X1 _3922_ (.A1(_0834_),
    .A2(net86),
    .A3(net81),
    .A4(_0835_),
    .ZN(_0969_));
 NAND2_X1 _3923_ (.A1(_0968_),
    .A2(_0969_),
    .ZN(_0970_));
 NAND2_X1 _3924_ (.A1(_0970_),
    .A2(net83),
    .ZN(_0971_));
 NAND3_X1 _3925_ (.A1(_0845_),
    .A2(_0846_),
    .A3(net85),
    .ZN(_0972_));
 NAND3_X1 _3926_ (.A1(_0838_),
    .A2(_0305_),
    .A3(_0839_),
    .ZN(_0973_));
 NAND3_X1 _3927_ (.A1(_0972_),
    .A2(_0973_),
    .A3(_0565_),
    .ZN(_0974_));
 NAND2_X1 _3928_ (.A1(_0971_),
    .A2(_0974_),
    .ZN(_0975_));
 NAND2_X1 _3929_ (.A1(_0975_),
    .A2(_0447_),
    .ZN(_0976_));
 NOR2_X1 _3930_ (.A1(_0575_),
    .A2(_0976_),
    .ZN(_0977_));
 AND3_X1 _3931_ (.A1(_2155_),
    .A2(_0967_),
    .A3(_0977_),
    .ZN(_0978_));
 NAND2_X2 _3932_ (.A1(_0944_),
    .A2(_0978_),
    .ZN(_0979_));
 AOI21_X1 _3933_ (.A(_0344_),
    .B1(_0563_),
    .B2(_0564_),
    .ZN(_0980_));
 AOI21_X1 _3934_ (.A(net84),
    .B1(_0559_),
    .B2(_0305_),
    .ZN(_0981_));
 OAI21_X1 _3935_ (.A(_0424_),
    .B1(_0980_),
    .B2(_0981_),
    .ZN(_0982_));
 NAND3_X1 _3936_ (.A1(_0501_),
    .A2(net115),
    .A3(_0502_),
    .ZN(_0983_));
 OAI21_X1 _3937_ (.A(net81),
    .B1(_0983_),
    .B2(net84),
    .ZN(_0984_));
 AND3_X1 _3938_ (.A1(_0982_),
    .A2(_0447_),
    .A3(_0984_),
    .ZN(_2191_));
 NAND2_X1 _3939_ (.A1(_0964_),
    .A2(_0344_),
    .ZN(_0985_));
 NAND3_X1 _3940_ (.A1(_0899_),
    .A2(_0344_),
    .A3(net87),
    .ZN(_0986_));
 AOI21_X1 _3941_ (.A(_0317_),
    .B1(_0986_),
    .B2(net81),
    .ZN(_0987_));
 NAND2_X1 _3942_ (.A1(_0960_),
    .A2(net83),
    .ZN(_0988_));
 NAND3_X1 _3943_ (.A1(_0985_),
    .A2(_0987_),
    .A3(_0988_),
    .ZN(_0989_));
 INV_X1 _3944_ (.A(_0989_),
    .ZN(_0990_));
 NAND2_X1 _3945_ (.A1(_2191_),
    .A2(_0990_),
    .ZN(_0991_));
 NAND2_X1 _3946_ (.A1(_0851_),
    .A2(_0305_),
    .ZN(_0992_));
 AOI21_X1 _3947_ (.A(_0317_),
    .B1(_0992_),
    .B2(_0341_),
    .ZN(_0993_));
 NAND3_X1 _3948_ (.A1(_0834_),
    .A2(net86),
    .A3(_0835_),
    .ZN(_0994_));
 OAI21_X1 _3949_ (.A(net81),
    .B1(_0994_),
    .B2(net83),
    .ZN(_0995_));
 NAND2_X1 _3950_ (.A1(_0993_),
    .A2(_0995_),
    .ZN(_0996_));
 AOI21_X1 _3951_ (.A(_0344_),
    .B1(_0973_),
    .B2(_0972_),
    .ZN(_0997_));
 NOR2_X1 _3952_ (.A1(_0996_),
    .A2(_0997_),
    .ZN(_0998_));
 NAND2_X1 _3953_ (.A1(_2187_),
    .A2(_0998_),
    .ZN(_0999_));
 NOR2_X1 _3954_ (.A1(_0991_),
    .A2(_0999_),
    .ZN(_1000_));
 OAI21_X1 _3955_ (.A(_0469_),
    .B1(_2120_),
    .B2(_0580_),
    .ZN(_1001_));
 AOI21_X1 _3956_ (.A(_0445_),
    .B1(_1001_),
    .B2(_0424_),
    .ZN(_1002_));
 AND3_X1 _3957_ (.A1(_1002_),
    .A2(_0316_),
    .A3(_0315_),
    .ZN(_1003_));
 AOI21_X1 _3958_ (.A(_0424_),
    .B1(_0657_),
    .B2(_0344_),
    .ZN(_1004_));
 NAND2_X1 _3959_ (.A1(_0630_),
    .A2(net82),
    .ZN(_1005_));
 AOI21_X1 _3960_ (.A(_0317_),
    .B1(_0587_),
    .B2(_0341_),
    .ZN(_1006_));
 NAND2_X1 _3961_ (.A1(_1005_),
    .A2(_1006_),
    .ZN(_1007_));
 NOR2_X1 _3962_ (.A1(_1004_),
    .A2(_1007_),
    .ZN(_1008_));
 NAND2_X1 _3963_ (.A1(_2179_),
    .A2(_1008_),
    .ZN(_1009_));
 INV_X1 _3964_ (.A(_1009_),
    .ZN(_1010_));
 AOI21_X1 _3965_ (.A(_0317_),
    .B1(_0948_),
    .B2(_0341_),
    .ZN(_1011_));
 AND3_X1 _3966_ (.A1(_0946_),
    .A2(_0344_),
    .A3(net86),
    .ZN(_1012_));
 OAI21_X1 _3967_ (.A(_1011_),
    .B1(_1012_),
    .B2(_0424_),
    .ZN(_1013_));
 NOR2_X1 _3968_ (.A1(_0954_),
    .A2(_0344_),
    .ZN(_1014_));
 NOR2_X1 _3969_ (.A1(_1013_),
    .A2(_1014_),
    .ZN(_1015_));
 NAND4_X2 _3970_ (.A1(_1000_),
    .A2(_1003_),
    .A3(_1010_),
    .A4(_1015_),
    .ZN(_1016_));
 NOR2_X4 _3971_ (.A1(_1016_),
    .A2(_0979_),
    .ZN(_1017_));
 NAND2_X4 _3972_ (.A1(net147),
    .A2(_1017_),
    .ZN(_1018_));
 NAND2_X1 _3973_ (.A1(_0906_),
    .A2(_1018_),
    .ZN(_1019_));
 TAPCELL_X1 PHY_16 ();
 TAPCELL_X1 PHY_15 ();
 NAND3_X1 _3976_ (.A1(_1017_),
    .A2(_2151_),
    .A3(net147),
    .ZN(_1022_));
 NAND2_X1 _3977_ (.A1(_1019_),
    .A2(_1022_),
    .ZN(net49));
 TAPCELL_X1 PHY_14 ();
 NAND2_X1 _3979_ (.A1(_1018_),
    .A2(_2151_),
    .ZN(_1024_));
 NAND3_X1 _3980_ (.A1(_1017_),
    .A2(_2154_),
    .A3(net147),
    .ZN(_1025_));
 NAND2_X1 _3981_ (.A1(_1024_),
    .A2(_1025_),
    .ZN(net60));
 NAND2_X1 _3982_ (.A1(net192),
    .A2(_2154_),
    .ZN(_1026_));
 XNOR2_X1 _3983_ (.A(_0957_),
    .B(_2153_),
    .ZN(_1027_));
 NAND3_X1 _3984_ (.A1(_1017_),
    .A2(net147),
    .A3(_1027_),
    .ZN(_1028_));
 NAND2_X1 _3985_ (.A1(_1026_),
    .A2(_1028_),
    .ZN(net71));
 NAND2_X1 _3986_ (.A1(_1018_),
    .A2(_1027_),
    .ZN(_1029_));
 NAND3_X1 _3987_ (.A1(_1017_),
    .A2(_2158_),
    .A3(net147),
    .ZN(_1030_));
 NAND2_X1 _3988_ (.A1(_1029_),
    .A2(_1030_),
    .ZN(net74));
 NAND2_X1 _3989_ (.A1(net193),
    .A2(_2158_),
    .ZN(_1031_));
 XNOR2_X1 _3990_ (.A(_0976_),
    .B(_2157_),
    .ZN(_1032_));
 NAND3_X1 _3991_ (.A1(_1017_),
    .A2(net147),
    .A3(_1032_),
    .ZN(_1033_));
 NAND2_X1 _3992_ (.A1(_1031_),
    .A2(_1033_),
    .ZN(net75));
 AND2_X1 _3993_ (.A1(_2155_),
    .A2(_0977_),
    .ZN(_2160_));
 NAND2_X1 _3994_ (.A1(net192),
    .A2(_1032_),
    .ZN(_1034_));
 NAND3_X1 _3995_ (.A1(net187),
    .A2(_2162_),
    .A3(net127),
    .ZN(_1035_));
 NAND2_X1 _3996_ (.A1(_1034_),
    .A2(_1035_),
    .ZN(net76));
 NAND2_X1 _3997_ (.A1(net192),
    .A2(_2162_),
    .ZN(_1036_));
 XNOR2_X1 _3998_ (.A(_0966_),
    .B(_2161_),
    .ZN(_1037_));
 NAND3_X1 _3999_ (.A1(net187),
    .A2(net127),
    .A3(_1037_),
    .ZN(_1038_));
 NAND2_X1 _4000_ (.A1(_1036_),
    .A2(_1038_),
    .ZN(net77));
 NAND2_X1 _4001_ (.A1(net192),
    .A2(_1037_),
    .ZN(_1039_));
 NAND3_X1 _4002_ (.A1(net187),
    .A2(_2166_),
    .A3(net147),
    .ZN(_1040_));
 NAND2_X1 _4003_ (.A1(_1039_),
    .A2(_1040_),
    .ZN(net78));
 NAND2_X1 _4004_ (.A1(net192),
    .A2(_2166_),
    .ZN(_1041_));
 XNOR2_X1 _4005_ (.A(_0941_),
    .B(_2165_),
    .ZN(_1042_));
 NAND3_X1 _4006_ (.A1(net187),
    .A2(net127),
    .A3(_1042_),
    .ZN(_1043_));
 NAND2_X1 _4007_ (.A1(_1041_),
    .A2(_1043_),
    .ZN(net79));
 NAND4_X4 _4008_ (.A1(_2155_),
    .A2(_0942_),
    .A3(_0967_),
    .A4(_0977_),
    .ZN(_1044_));
 INV_X1 _4009_ (.A(_1044_),
    .ZN(_2168_));
 NAND2_X1 _4010_ (.A1(net192),
    .A2(_1042_),
    .ZN(_1045_));
 NAND3_X1 _4011_ (.A1(net187),
    .A2(_2170_),
    .A3(net147),
    .ZN(_1046_));
 NAND2_X1 _4012_ (.A1(_1045_),
    .A2(_1046_),
    .ZN(net80));
 NAND2_X1 _4013_ (.A1(net193),
    .A2(_2170_),
    .ZN(_1047_));
 TAPCELL_X1 PHY_13 ();
 XNOR2_X1 _4015_ (.A(_0929_),
    .B(_2169_),
    .ZN(_1049_));
 NAND3_X1 _4016_ (.A1(net187),
    .A2(net127),
    .A3(_1049_),
    .ZN(_1050_));
 NAND2_X1 _4017_ (.A1(_1047_),
    .A2(_1050_),
    .ZN(net50));
 TAPCELL_X1 PHY_12 ();
 NAND2_X1 _4019_ (.A1(net192),
    .A2(_1049_),
    .ZN(_1052_));
 NAND3_X1 _4020_ (.A1(net182),
    .A2(_2174_),
    .A3(net127),
    .ZN(_1053_));
 NAND2_X1 _4021_ (.A1(_1052_),
    .A2(_1053_),
    .ZN(net51));
 NAND2_X1 _4022_ (.A1(net192),
    .A2(_2174_),
    .ZN(_1054_));
 XNOR2_X1 _4023_ (.A(_0912_),
    .B(_2173_),
    .ZN(_1055_));
 NAND3_X1 _4024_ (.A1(net182),
    .A2(net127),
    .A3(_1055_),
    .ZN(_1056_));
 NAND2_X1 _4025_ (.A1(_1054_),
    .A2(_1056_),
    .ZN(net52));
 NOR2_X4 _4026_ (.A1(_0930_),
    .A2(_1044_),
    .ZN(_2171_));
 AND2_X1 _4027_ (.A1(_0913_),
    .A2(_2171_),
    .ZN(_2175_));
 NAND2_X1 _4028_ (.A1(net192),
    .A2(_1055_),
    .ZN(_1057_));
 NAND3_X1 _4029_ (.A1(net182),
    .A2(_2178_),
    .A3(net127),
    .ZN(_1058_));
 NAND2_X1 _4030_ (.A1(_1057_),
    .A2(_1058_),
    .ZN(net53));
 NAND2_X1 _4031_ (.A1(net192),
    .A2(_2178_),
    .ZN(_1059_));
 XNOR2_X1 _4032_ (.A(_2177_),
    .B(_0908_),
    .ZN(_1060_));
 NAND3_X1 _4033_ (.A1(net182),
    .A2(net127),
    .A3(_1060_),
    .ZN(_1061_));
 NAND2_X1 _4034_ (.A1(_1059_),
    .A2(_1061_),
    .ZN(net54));
 NAND2_X1 _4035_ (.A1(net193),
    .A2(_1060_),
    .ZN(_1062_));
 NAND3_X1 _4036_ (.A1(net182),
    .A2(_2182_),
    .A3(net127),
    .ZN(_1063_));
 NAND2_X1 _4037_ (.A1(_1062_),
    .A2(_1063_),
    .ZN(net55));
 NAND2_X1 _4038_ (.A1(net192),
    .A2(_2182_),
    .ZN(_1064_));
 XOR2_X1 _4039_ (.A(_1008_),
    .B(_2181_),
    .Z(_1065_));
 NAND3_X1 _4040_ (.A1(net182),
    .A2(_1065_),
    .A3(net127),
    .ZN(_1066_));
 NAND2_X1 _4041_ (.A1(_1064_),
    .A2(_1066_),
    .ZN(net56));
 NAND3_X4 _4042_ (.A1(_2171_),
    .A2(_0909_),
    .A3(_0913_),
    .ZN(_1067_));
 NOR2_X4 _4043_ (.A1(_1009_),
    .A2(_1067_),
    .ZN(_2184_));
 NAND2_X1 _4044_ (.A1(net193),
    .A2(_1065_),
    .ZN(_1068_));
 NAND3_X1 _4045_ (.A1(net182),
    .A2(_2186_),
    .A3(net127),
    .ZN(_1069_));
 NAND2_X1 _4046_ (.A1(_1068_),
    .A2(_1069_),
    .ZN(net57));
 NAND2_X1 _4047_ (.A1(_1018_),
    .A2(_2186_),
    .ZN(_1070_));
 INV_X1 _4048_ (.A(_1015_),
    .ZN(_1071_));
 XNOR2_X2 _4049_ (.A(_1071_),
    .B(_2185_),
    .ZN(_1072_));
 NAND3_X1 _4050_ (.A1(net182),
    .A2(net127),
    .A3(_1072_),
    .ZN(_1073_));
 NAND2_X1 _4051_ (.A1(_1073_),
    .A2(_1070_),
    .ZN(net58));
 NAND2_X1 _4052_ (.A1(_1018_),
    .A2(_1072_),
    .ZN(_1074_));
 NAND3_X1 _4053_ (.A1(net182),
    .A2(_2190_),
    .A3(net127),
    .ZN(_1075_));
 NAND2_X1 _4054_ (.A1(_1075_),
    .A2(_1074_),
    .ZN(net59));
 NAND2_X1 _4055_ (.A1(_1018_),
    .A2(_2190_),
    .ZN(_1076_));
 XOR2_X1 _4056_ (.A(_2189_),
    .B(_0998_),
    .Z(_1077_));
 NAND3_X1 _4057_ (.A1(net182),
    .A2(net127),
    .A3(_1077_),
    .ZN(_1078_));
 NAND2_X1 _4058_ (.A1(_1078_),
    .A2(_1076_),
    .ZN(net61));
 INV_X1 _4059_ (.A(_0999_),
    .ZN(_1079_));
 NOR2_X1 _4060_ (.A1(_0476_),
    .A2(_1071_),
    .ZN(_1080_));
 NAND3_X4 _4061_ (.A1(_2184_),
    .A2(_1079_),
    .A3(_1080_),
    .ZN(_1081_));
 INV_X1 _4062_ (.A(_1081_),
    .ZN(_2192_));
 NAND2_X1 _4063_ (.A1(net193),
    .A2(_1077_),
    .ZN(_1082_));
 NAND3_X1 _4064_ (.A1(net182),
    .A2(_2194_),
    .A3(net127),
    .ZN(_1083_));
 NAND2_X1 _4065_ (.A1(_1082_),
    .A2(_1083_),
    .ZN(net62));
 NAND2_X1 _4066_ (.A1(net193),
    .A2(_2194_),
    .ZN(_1084_));
 XNOR2_X1 _4067_ (.A(_0989_),
    .B(_2193_),
    .ZN(_1085_));
 NAND3_X1 _4068_ (.A1(net182),
    .A2(net127),
    .A3(_1085_),
    .ZN(_1086_));
 NAND2_X1 _4069_ (.A1(_1084_),
    .A2(_1086_),
    .ZN(net63));
 INV_X1 _4070_ (.A(_2088_),
    .ZN(_2109_));
 NOR4_X1 _4071_ (.A1(_2073_),
    .A2(_2081_),
    .A3(_0211_),
    .A4(_2109_),
    .ZN(_1087_));
 NOR2_X1 _4072_ (.A1(net118),
    .A2(_2267_),
    .ZN(_1088_));
 INV_X1 _4073_ (.A(_2270_),
    .ZN(_2268_));
 TAPCELL_X1 PHY_11 ();
 AOI21_X1 _4075_ (.A(_1088_),
    .B1(_2268_),
    .B2(net118),
    .ZN(_1090_));
 NAND4_X1 _4076_ (.A1(_1087_),
    .A2(_2069_),
    .A3(_2139_),
    .A4(_1090_),
    .ZN(_1091_));
 NOR2_X1 _4077_ (.A1(_1091_),
    .A2(_1975_),
    .ZN(_2042_));
 INV_X1 _4078_ (.A(_2074_),
    .ZN(_2057_));
 INV_X1 _4079_ (.A(_2050_),
    .ZN(net65));
 INV_X1 _4080_ (.A(_2054_),
    .ZN(net66));
 INV_X1 _4081_ (.A(_2063_),
    .ZN(net70));
 INV_X1 _4082_ (.A(_2076_),
    .ZN(_2072_));
 NOR2_X1 _4083_ (.A1(_1091_),
    .A2(_0210_),
    .ZN(_2106_));
 NAND2_X2 _4084_ (.A1(_0229_),
    .A2(_2072_),
    .ZN(_1092_));
 XNOR2_X1 _4085_ (.A(_2077_),
    .B(_2097_),
    .ZN(_1093_));
 OAI21_X4 _4086_ (.A(_1092_),
    .B1(_1093_),
    .B2(_0229_),
    .ZN(_2111_));
 INV_X1 _4087_ (.A(_0241_),
    .ZN(_2121_));
 INV_X1 _4088_ (.A(_2129_),
    .ZN(_2125_));
 INV_X1 _4089_ (.A(_2090_),
    .ZN(_2047_));
 NOR2_X4 _4090_ (.A1(_0867_),
    .A2(_0902_),
    .ZN(_2148_));
 NAND2_X1 _4091_ (.A1(_2160_),
    .A2(_0967_),
    .ZN(_1094_));
 INV_X1 _4092_ (.A(_1094_),
    .ZN(_2163_));
 NAND2_X1 _4093_ (.A1(_2240_),
    .A2(net90),
    .ZN(_1095_));
 OAI21_X1 _4094_ (.A(_1095_),
    .B1(net31),
    .B2(net90),
    .ZN(_1096_));
 XNOR2_X1 _4095_ (.A(_1648_),
    .B(_1096_),
    .ZN(_1097_));
 INV_X1 _4096_ (.A(_1097_),
    .ZN(_2272_));
 NAND2_X1 _4097_ (.A1(_2243_),
    .A2(net90),
    .ZN(_1098_));
 OAI21_X1 _4098_ (.A(_1098_),
    .B1(net30),
    .B2(net90),
    .ZN(_1099_));
 XNOR2_X1 _4099_ (.A(_1648_),
    .B(_1099_),
    .ZN(_1100_));
 INV_X1 _4100_ (.A(_1100_),
    .ZN(_1977_));
 TAPCELL_X1 PHY_10 ();
 NOR2_X1 _4102_ (.A1(net90),
    .A2(net29),
    .ZN(_1102_));
 AOI21_X1 _4103_ (.A(_1102_),
    .B1(_2246_),
    .B2(net90),
    .ZN(_1103_));
 XNOR2_X1 _4104_ (.A(_1648_),
    .B(_1103_),
    .ZN(_2278_));
 NOR2_X1 _4105_ (.A1(net90),
    .A2(net27),
    .ZN(_1104_));
 AOI21_X1 _4106_ (.A(_1104_),
    .B1(_2249_),
    .B2(net90),
    .ZN(_1105_));
 XNOR2_X2 _4107_ (.A(_1648_),
    .B(_1105_),
    .ZN(_1982_));
 TAPCELL_X1 PHY_9 ();
 NAND2_X1 _4109_ (.A1(_1783_),
    .A2(net95),
    .ZN(_1107_));
 OAI21_X1 _4110_ (.A(_1107_),
    .B1(net95),
    .B2(_1801_),
    .ZN(_1108_));
 NAND2_X1 _4111_ (.A1(_1108_),
    .A2(net129),
    .ZN(_1109_));
 OAI21_X1 _4112_ (.A(_1617_),
    .B1(_1777_),
    .B2(_1570_),
    .ZN(_1110_));
 OAI21_X1 _4113_ (.A(_1110_),
    .B1(_1771_),
    .B2(_1617_),
    .ZN(_1111_));
 NAND2_X1 _4114_ (.A1(_1111_),
    .A2(_1546_),
    .ZN(_1112_));
 NAND2_X1 _4115_ (.A1(_1109_),
    .A2(_1112_),
    .ZN(_1113_));
 NAND2_X1 _4116_ (.A1(_1113_),
    .A2(net105),
    .ZN(_1114_));
 NOR3_X1 _4117_ (.A1(_1570_),
    .A2(net95),
    .A3(_1633_),
    .ZN(_1115_));
 INV_X1 _4118_ (.A(_1793_),
    .ZN(_1116_));
 AOI21_X1 _4119_ (.A(_1115_),
    .B1(_1116_),
    .B2(net95),
    .ZN(_1117_));
 NOR2_X1 _4120_ (.A1(_1117_),
    .A2(net129),
    .ZN(_1118_));
 INV_X1 _4121_ (.A(_1118_),
    .ZN(_1119_));
 NAND2_X1 _4122_ (.A1(_1119_),
    .A2(_1576_),
    .ZN(_1120_));
 NAND2_X1 _4123_ (.A1(_1114_),
    .A2(_1120_),
    .ZN(_1121_));
 NOR3_X1 _4124_ (.A1(_1121_),
    .A2(_1814_),
    .A3(_1643_),
    .ZN(_1122_));
 XNOR2_X1 _4125_ (.A(_1627_),
    .B(_1122_),
    .ZN(_2284_));
 NAND3_X1 _4126_ (.A1(_1836_),
    .A2(_1565_),
    .A3(net98),
    .ZN(_1123_));
 XNOR2_X1 _4127_ (.A(_1627_),
    .B(_1123_),
    .ZN(_1124_));
 INV_X1 _4128_ (.A(_1124_),
    .ZN(_1987_));
 NOR2_X1 _4129_ (.A1(net90),
    .A2(net24),
    .ZN(_1125_));
 AOI21_X1 _4130_ (.A(_1125_),
    .B1(_2258_),
    .B2(net90),
    .ZN(_1126_));
 XNOR2_X1 _4131_ (.A(_1648_),
    .B(_1126_),
    .ZN(_2290_));
 NOR2_X1 _4132_ (.A1(net90),
    .A2(net23),
    .ZN(_1127_));
 AOI21_X2 _4133_ (.A(_1127_),
    .B1(_2261_),
    .B2(net90),
    .ZN(_1128_));
 XNOR2_X2 _4134_ (.A(_1648_),
    .B(_1128_),
    .ZN(_1992_));
 NOR2_X1 _4135_ (.A1(net90),
    .A2(net22),
    .ZN(_1129_));
 AOI21_X1 _4136_ (.A(_1129_),
    .B1(_2264_),
    .B2(net90),
    .ZN(_1130_));
 XNOR2_X1 _4137_ (.A(_1648_),
    .B(_1130_),
    .ZN(_2296_));
 INV_X1 _4138_ (.A(_1997_),
    .ZN(_2300_));
 OR2_X1 _4139_ (.A1(_1108_),
    .A2(net129),
    .ZN(_1131_));
 OR2_X1 _4140_ (.A1(_1117_),
    .A2(net110),
    .ZN(_1132_));
 NAND2_X1 _4141_ (.A1(_1131_),
    .A2(_1132_),
    .ZN(_1133_));
 NAND2_X1 _4142_ (.A1(_1133_),
    .A2(net105),
    .ZN(_1134_));
 NAND2_X1 _4143_ (.A1(_1134_),
    .A2(_1643_),
    .ZN(_1135_));
 NAND2_X1 _4144_ (.A1(_1111_),
    .A2(net129),
    .ZN(_1136_));
 NAND2_X1 _4145_ (.A1(_1765_),
    .A2(_1617_),
    .ZN(_1137_));
 OAI21_X1 _4146_ (.A(_1137_),
    .B1(_1617_),
    .B2(_1757_),
    .ZN(_1138_));
 NAND2_X1 _4147_ (.A1(_1138_),
    .A2(net110),
    .ZN(_1139_));
 NAND3_X1 _4148_ (.A1(_1136_),
    .A2(_1576_),
    .A3(_1139_),
    .ZN(_1140_));
 NOR2_X1 _4149_ (.A1(_1825_),
    .A2(_1617_),
    .ZN(_1141_));
 AOI21_X1 _4150_ (.A(_1141_),
    .B1(_1744_),
    .B2(_1617_),
    .ZN(_1142_));
 NAND2_X1 _4151_ (.A1(_1737_),
    .A2(net94),
    .ZN(_1143_));
 INV_X1 _4152_ (.A(_1750_),
    .ZN(_1144_));
 OAI21_X1 _4153_ (.A(_1143_),
    .B1(_1144_),
    .B2(net94),
    .ZN(_1145_));
 MUX2_X1 _4154_ (.A(_1142_),
    .B(_1145_),
    .S(_1620_),
    .Z(_1146_));
 INV_X1 _4155_ (.A(_1146_),
    .ZN(_1147_));
 NAND2_X1 _4156_ (.A1(_1147_),
    .A2(net105),
    .ZN(_1148_));
 NAND3_X1 _4157_ (.A1(_1140_),
    .A2(net89),
    .A3(_1148_),
    .ZN(_1149_));
 NAND3_X1 _4158_ (.A1(_1135_),
    .A2(_1149_),
    .A3(_1565_),
    .ZN(_1150_));
 XNOR2_X1 _4159_ (.A(_1627_),
    .B(_1150_),
    .ZN(_1151_));
 INV_X1 _4160_ (.A(_1151_),
    .ZN(_2304_));
 NOR2_X1 _4161_ (.A1(net90),
    .A2(_1826_),
    .ZN(_1152_));
 XNOR2_X2 _4162_ (.A(_1648_),
    .B(_1152_),
    .ZN(_2002_));
 NOR2_X1 _4163_ (.A1(net90),
    .A2(_1815_),
    .ZN(_1153_));
 XNOR2_X1 _4164_ (.A(_1648_),
    .B(_1153_),
    .ZN(_2310_));
 INV_X1 _4165_ (.A(_2007_),
    .ZN(_2314_));
 NOR2_X1 _4166_ (.A1(net90),
    .A2(_1854_),
    .ZN(_1154_));
 XNOR2_X1 _4167_ (.A(_1648_),
    .B(_1154_),
    .ZN(_2318_));
 INV_X1 _4168_ (.A(_2012_),
    .ZN(_2322_));
 NAND3_X1 _4169_ (.A1(_1109_),
    .A2(_1576_),
    .A3(_1112_),
    .ZN(_1155_));
 MUX2_X1 _4170_ (.A(_1145_),
    .B(_1138_),
    .S(_1620_),
    .Z(_1156_));
 OR2_X1 _4171_ (.A1(_1156_),
    .A2(_1576_),
    .ZN(_1157_));
 NAND3_X1 _4172_ (.A1(_1155_),
    .A2(_1157_),
    .A3(_1643_),
    .ZN(_1158_));
 OAI21_X1 _4173_ (.A(net93),
    .B1(_1570_),
    .B2(_1817_),
    .ZN(_1159_));
 INV_X1 _4174_ (.A(_1828_),
    .ZN(_1160_));
 OAI21_X1 _4175_ (.A(_1159_),
    .B1(_1160_),
    .B2(net93),
    .ZN(_1161_));
 MUX2_X1 _4176_ (.A(_1161_),
    .B(_1142_),
    .S(net145),
    .Z(_1162_));
 NAND2_X1 _4177_ (.A1(_1162_),
    .A2(_1576_),
    .ZN(_1163_));
 NAND2_X1 _4178_ (.A1(_1856_),
    .A2(net93),
    .ZN(_1164_));
 OAI21_X1 _4179_ (.A(_1164_),
    .B1(_1821_),
    .B2(net93),
    .ZN(_1165_));
 INV_X1 _4180_ (.A(_1165_),
    .ZN(_1166_));
 NAND2_X1 _4181_ (.A1(_1166_),
    .A2(net145),
    .ZN(_1167_));
 OAI21_X1 _4182_ (.A(net93),
    .B1(_1570_),
    .B2(_1872_),
    .ZN(_1168_));
 INV_X1 _4183_ (.A(_1858_),
    .ZN(_1169_));
 OAI21_X1 _4184_ (.A(_1168_),
    .B1(net93),
    .B2(_1169_),
    .ZN(_1170_));
 OAI21_X1 _4185_ (.A(_1167_),
    .B1(net129),
    .B2(_1170_),
    .ZN(_1171_));
 OAI21_X1 _4186_ (.A(_1163_),
    .B1(_1576_),
    .B2(_1171_),
    .ZN(_1172_));
 AOI21_X1 _4187_ (.A(_1814_),
    .B1(_1172_),
    .B2(net89),
    .ZN(_1173_));
 NOR2_X1 _4188_ (.A1(_1119_),
    .A2(_1576_),
    .ZN(_1174_));
 INV_X1 _4189_ (.A(_1174_),
    .ZN(_1175_));
 NOR2_X1 _4190_ (.A1(_1175_),
    .A2(_1643_),
    .ZN(_1176_));
 AOI22_X1 _4191_ (.A1(_1158_),
    .A2(_1173_),
    .B1(_1176_),
    .B2(_1843_),
    .ZN(_1177_));
 XNOR2_X1 _4192_ (.A(_1177_),
    .B(_1627_),
    .ZN(_1178_));
 INV_X1 _4193_ (.A(_1178_),
    .ZN(_2326_));
 INV_X1 _4194_ (.A(_2017_),
    .ZN(_2330_));
 NOR2_X1 _4195_ (.A1(net90),
    .A2(_1900_),
    .ZN(_1179_));
 XNOR2_X1 _4196_ (.A(_1648_),
    .B(_1179_),
    .ZN(_2334_));
 INV_X1 _4197_ (.A(_2021_),
    .ZN(_2338_));
 MUX2_X1 _4198_ (.A(_1162_),
    .B(_1156_),
    .S(_1576_),
    .Z(_1180_));
 NAND2_X1 _4199_ (.A1(_1180_),
    .A2(_1643_),
    .ZN(_1181_));
 OAI21_X1 _4200_ (.A(_1617_),
    .B1(_1570_),
    .B2(_1876_),
    .ZN(_1182_));
 OAI21_X1 _4201_ (.A(_1182_),
    .B1(_1902_),
    .B2(_1617_),
    .ZN(_1183_));
 NAND2_X1 _4202_ (.A1(_1183_),
    .A2(net129),
    .ZN(_1184_));
 NAND2_X1 _4203_ (.A1(_1906_),
    .A2(_1617_),
    .ZN(_1185_));
 OAI21_X1 _4204_ (.A(_1185_),
    .B1(_1617_),
    .B2(_1921_),
    .ZN(_1186_));
 INV_X1 _4205_ (.A(_1186_),
    .ZN(_1187_));
 OAI21_X1 _4206_ (.A(_1184_),
    .B1(_1187_),
    .B2(net145),
    .ZN(_1188_));
 NAND2_X1 _4207_ (.A1(_1188_),
    .A2(net111),
    .ZN(_1189_));
 OAI21_X1 _4208_ (.A(_1189_),
    .B1(_1171_),
    .B2(net105),
    .ZN(_1190_));
 AOI21_X1 _4209_ (.A(_1814_),
    .B1(_1190_),
    .B2(net89),
    .ZN(_1191_));
 NAND2_X1 _4210_ (.A1(_1181_),
    .A2(_1191_),
    .ZN(_1192_));
 NAND3_X1 _4211_ (.A1(_1114_),
    .A2(net89),
    .A3(_1120_),
    .ZN(_1193_));
 OAI21_X1 _4212_ (.A(_1192_),
    .B1(_1884_),
    .B2(_1193_),
    .ZN(_1194_));
 TAPCELL_X1 PHY_8 ();
 XNOR2_X1 _4214_ (.A(_1194_),
    .B(_1733_),
    .ZN(_1196_));
 INV_X1 _4215_ (.A(_1196_),
    .ZN(_2342_));
 INV_X1 _4216_ (.A(_2026_),
    .ZN(_2346_));
 OR2_X1 _4217_ (.A1(_1183_),
    .A2(net145),
    .ZN(_1197_));
 OAI21_X1 _4218_ (.A(_1197_),
    .B1(net102),
    .B2(_1170_),
    .ZN(_1198_));
 INV_X1 _4219_ (.A(net17),
    .ZN(_1199_));
 NOR2_X1 _4220_ (.A1(net109),
    .A2(_1199_),
    .ZN(_1200_));
 NAND2_X1 _4221_ (.A1(_1571_),
    .A2(_1200_),
    .ZN(_1201_));
 MUX2_X1 _4222_ (.A(_1201_),
    .B(_1925_),
    .S(_1617_),
    .Z(_1202_));
 OAI21_X1 _4223_ (.A(_1553_),
    .B1(_1202_),
    .B2(net129),
    .ZN(_1203_));
 NOR2_X1 _4224_ (.A1(_1186_),
    .A2(net102),
    .ZN(_1204_));
 OAI22_X1 _4225_ (.A1(_1198_),
    .A2(net105),
    .B1(_1203_),
    .B2(_1204_),
    .ZN(_1205_));
 AOI21_X1 _4226_ (.A(_1814_),
    .B1(_1205_),
    .B2(net89),
    .ZN(_1206_));
 NAND2_X1 _4227_ (.A1(_1161_),
    .A2(net129),
    .ZN(_1207_));
 OAI21_X1 _4228_ (.A(_1207_),
    .B1(_1166_),
    .B2(net145),
    .ZN(_1208_));
 NOR2_X1 _4229_ (.A1(_1208_),
    .A2(_1576_),
    .ZN(_1209_));
 AOI21_X1 _4230_ (.A(_1209_),
    .B1(_1147_),
    .B2(_1576_),
    .ZN(_1210_));
 INV_X1 _4231_ (.A(_1210_),
    .ZN(_1211_));
 OAI21_X1 _4232_ (.A(_1206_),
    .B1(_1211_),
    .B2(net89),
    .ZN(_1212_));
 NAND3_X1 _4233_ (.A1(_1131_),
    .A2(_1132_),
    .A3(_1576_),
    .ZN(_1213_));
 NAND2_X1 _4234_ (.A1(_1136_),
    .A2(_1139_),
    .ZN(_1214_));
 NAND2_X1 _4235_ (.A1(_1214_),
    .A2(net111),
    .ZN(_1215_));
 NAND3_X1 _4236_ (.A1(_1213_),
    .A2(net89),
    .A3(_1215_),
    .ZN(_1216_));
 OAI21_X1 _4237_ (.A(_1212_),
    .B1(_1216_),
    .B2(_1884_),
    .ZN(_1217_));
 XNOR2_X1 _4238_ (.A(_1217_),
    .B(_1733_),
    .ZN(_1218_));
 INV_X1 _4239_ (.A(_1218_),
    .ZN(_2350_));
 NAND3_X1 _4240_ (.A1(_1847_),
    .A2(net97),
    .A3(_1851_),
    .ZN(_1219_));
 NAND2_X1 _4241_ (.A1(_1641_),
    .A2(_1643_),
    .ZN(_1220_));
 AND2_X1 _4242_ (.A1(_1219_),
    .A2(_1220_),
    .ZN(_1221_));
 NAND2_X1 _4243_ (.A1(_1221_),
    .A2(_1843_),
    .ZN(_1222_));
 AOI21_X1 _4244_ (.A(_1814_),
    .B1(_1862_),
    .B2(_1643_),
    .ZN(_1223_));
 AND2_X1 _4245_ (.A1(_1909_),
    .A2(_1576_),
    .ZN(_1224_));
 OAI21_X1 _4246_ (.A(net103),
    .B1(_1201_),
    .B2(net93),
    .ZN(_1225_));
 OAI21_X1 _4247_ (.A(_1225_),
    .B1(_1926_),
    .B2(net103),
    .ZN(_1226_));
 OAI21_X1 _4248_ (.A(net89),
    .B1(_1226_),
    .B2(_1576_),
    .ZN(_1227_));
 OAI21_X1 _4249_ (.A(_1223_),
    .B1(_1224_),
    .B2(_1227_),
    .ZN(_1228_));
 NAND2_X1 _4250_ (.A1(_1222_),
    .A2(_1228_),
    .ZN(_1229_));
 XNOR2_X1 _4251_ (.A(_1229_),
    .B(_1733_),
    .ZN(_1230_));
 INV_X1 _4252_ (.A(_1230_),
    .ZN(_2032_));
 NAND3_X1 _4253_ (.A1(_1155_),
    .A2(_1157_),
    .A3(net89),
    .ZN(_1231_));
 NAND2_X1 _4254_ (.A1(_1175_),
    .A2(_1643_),
    .ZN(_1232_));
 NAND3_X1 _4255_ (.A1(_1231_),
    .A2(_1843_),
    .A3(_1232_),
    .ZN(_1233_));
 NAND2_X1 _4256_ (.A1(_1172_),
    .A2(_1643_),
    .ZN(_1234_));
 NAND2_X1 _4257_ (.A1(net111),
    .A2(net129),
    .ZN(_1235_));
 OAI221_X1 _4258_ (.A(net89),
    .B1(_1202_),
    .B2(_1235_),
    .C1(_1188_),
    .C2(net111),
    .ZN(_1236_));
 NAND3_X1 _4259_ (.A1(_1234_),
    .A2(_1565_),
    .A3(_1236_),
    .ZN(_1237_));
 NAND2_X1 _4260_ (.A1(_1233_),
    .A2(_1237_),
    .ZN(_1238_));
 XNOR2_X1 _4261_ (.A(_1238_),
    .B(_1733_),
    .ZN(_1239_));
 INV_X1 _4262_ (.A(_1239_),
    .ZN(_2037_));
 AOI21_X4 _4263_ (.A(_1564_),
    .B1(_2373_),
    .B2(_2374_),
    .ZN(_2356_));
 XNOR2_X2 _4264_ (.A(_2358_),
    .B(_1569_),
    .ZN(_1240_));
 INV_X1 _4265_ (.A(_2359_),
    .ZN(_1241_));
 NAND2_X4 _4266_ (.A1(_1241_),
    .A2(_1240_),
    .ZN(_1242_));
 NOR3_X1 _4267_ (.A1(_1777_),
    .A2(net95),
    .A3(_1242_),
    .ZN(_1243_));
 INV_X8 _4268_ (.A(_1242_),
    .ZN(_1244_));
 TAPCELL_X1 PHY_7 ();
 TAPCELL_X1 PHY_6 ();
 NAND4_X1 _4271_ (.A1(_1775_),
    .A2(net95),
    .A3(_1776_),
    .A4(net128),
    .ZN(_1247_));
 NAND3_X1 _4272_ (.A1(_1764_),
    .A2(_1617_),
    .A3(net128),
    .ZN(_1248_));
 NAND2_X1 _4273_ (.A1(_1769_),
    .A2(net128),
    .ZN(_1249_));
 NAND3_X1 _4274_ (.A1(_1247_),
    .A2(_1248_),
    .A3(_1249_),
    .ZN(_1250_));
 TAPCELL_X1 PHY_5 ();
 INV_X2 _4276_ (.A(net88),
    .ZN(_1252_));
 TAPCELL_X1 PHY_4 ();
 AOI21_X1 _4278_ (.A(_1243_),
    .B1(_1250_),
    .B2(_1252_),
    .ZN(_1254_));
 OR2_X1 _4279_ (.A1(_1633_),
    .A2(_1252_),
    .ZN(_1255_));
 NAND2_X1 _4280_ (.A1(_1798_),
    .A2(_1255_),
    .ZN(_1256_));
 NAND2_X1 _4281_ (.A1(_1256_),
    .A2(net95),
    .ZN(_1257_));
 NAND2_X1 _4282_ (.A1(_1257_),
    .A2(_1781_),
    .ZN(_1258_));
 NAND2_X1 _4283_ (.A1(_1791_),
    .A2(_1792_),
    .ZN(_1259_));
 AOI21_X1 _4284_ (.A(_1252_),
    .B1(_1259_),
    .B2(_1798_),
    .ZN(_1260_));
 OAI21_X1 _4285_ (.A(net128),
    .B1(_1258_),
    .B2(_1260_),
    .ZN(_1261_));
 NAND2_X1 _4286_ (.A1(_1254_),
    .A2(_1261_),
    .ZN(_1262_));
 TAPCELL_X1 PHY_3 ();
 INV_X2 _4288_ (.A(_2372_),
    .ZN(_1264_));
 NAND2_X1 _4289_ (.A1(_1262_),
    .A2(_1264_),
    .ZN(_1265_));
 NAND3_X1 _4290_ (.A1(_1742_),
    .A2(_1617_),
    .A3(net128),
    .ZN(_1266_));
 NAND3_X1 _4291_ (.A1(_1734_),
    .A2(_1736_),
    .A3(net134),
    .ZN(_1267_));
 OAI21_X1 _4292_ (.A(_1266_),
    .B1(_1267_),
    .B2(_1617_),
    .ZN(_1268_));
 NAND2_X1 _4293_ (.A1(_1268_),
    .A2(_1252_),
    .ZN(_1269_));
 NAND2_X1 _4294_ (.A1(_1755_),
    .A2(net128),
    .ZN(_1270_));
 NAND2_X1 _4295_ (.A1(_1270_),
    .A2(net95),
    .ZN(_1271_));
 TAPCELL_X1 PHY_2 ();
 OAI21_X1 _4297_ (.A(_1617_),
    .B1(_1748_),
    .B2(_1242_),
    .ZN(_1273_));
 NAND3_X1 _4298_ (.A1(_1271_),
    .A2(_2363_),
    .A3(_1273_),
    .ZN(_1274_));
 NAND2_X1 _4299_ (.A1(_1269_),
    .A2(_1274_),
    .ZN(_1275_));
 NAND3_X1 _4300_ (.A1(_1742_),
    .A2(net94),
    .A3(net134),
    .ZN(_1276_));
 NAND2_X1 _4301_ (.A1(net134),
    .A2(_1824_),
    .ZN(_1277_));
 INV_X2 _4302_ (.A(_1277_),
    .ZN(_1278_));
 NAND2_X1 _4303_ (.A1(_1278_),
    .A2(_1617_),
    .ZN(_1279_));
 NAND2_X1 _4304_ (.A1(_1276_),
    .A2(_1279_),
    .ZN(_1280_));
 NAND2_X1 _4305_ (.A1(_1280_),
    .A2(_2363_),
    .ZN(_1281_));
 NAND2_X1 _4306_ (.A1(_1244_),
    .A2(_1827_),
    .ZN(_1282_));
 NAND2_X1 _4307_ (.A1(_1282_),
    .A2(net94),
    .ZN(_1283_));
 NOR2_X1 _4308_ (.A1(net135),
    .A2(_1817_),
    .ZN(_1284_));
 OAI21_X1 _4309_ (.A(_1283_),
    .B1(net94),
    .B2(_1284_),
    .ZN(_1285_));
 OAI21_X1 _4310_ (.A(_1281_),
    .B1(_2363_),
    .B2(_1285_),
    .ZN(_1286_));
 NOR2_X1 _4311_ (.A1(_1275_),
    .A2(_1286_),
    .ZN(_1287_));
 NAND2_X1 _4312_ (.A1(_1282_),
    .A2(_1617_),
    .ZN(_1288_));
 OAI21_X1 _4313_ (.A(_1288_),
    .B1(_1278_),
    .B2(_1617_),
    .ZN(_1289_));
 NAND4_X1 _4314_ (.A1(_1276_),
    .A2(_1252_),
    .A3(_1279_),
    .A4(_1289_),
    .ZN(_1290_));
 AND2_X1 _4315_ (.A1(_1734_),
    .A2(_1736_),
    .ZN(_1291_));
 NAND3_X1 _4316_ (.A1(_1291_),
    .A2(_1617_),
    .A3(net128),
    .ZN(_1292_));
 NAND3_X1 _4317_ (.A1(_1749_),
    .A2(net94),
    .A3(net128),
    .ZN(_1293_));
 NAND3_X1 _4318_ (.A1(_1292_),
    .A2(_1293_),
    .A3(_2363_),
    .ZN(_1294_));
 OAI21_X1 _4319_ (.A(_1290_),
    .B1(_1294_),
    .B2(_1268_),
    .ZN(_1295_));
 NAND2_X1 _4320_ (.A1(_1287_),
    .A2(_1295_),
    .ZN(_1296_));
 TAPCELL_X1 PHY_1 ();
 NAND2_X1 _4322_ (.A1(_1296_),
    .A2(_2372_),
    .ZN(_1298_));
 NAND2_X1 _4323_ (.A1(net134),
    .A2(_1200_),
    .ZN(_1299_));
 NOR3_X1 _4324_ (.A1(_1299_),
    .A2(_1617_),
    .A3(_1252_),
    .ZN(_1300_));
 AND2_X1 _4325_ (.A1(_1300_),
    .A2(_1264_),
    .ZN(_1301_));
 XNOR2_X1 _4326_ (.A(_1575_),
    .B(_2371_),
    .ZN(_1302_));
 INV_X2 _4327_ (.A(_1302_),
    .ZN(_1303_));
 NAND2_X1 _4328_ (.A1(_1301_),
    .A2(_1303_),
    .ZN(_1304_));
 INV_X1 _4329_ (.A(_2376_),
    .ZN(_1305_));
 NAND2_X1 _4330_ (.A1(_1304_),
    .A2(_1305_),
    .ZN(_1306_));
 NAND2_X1 _4331_ (.A1(_1244_),
    .A2(_1820_),
    .ZN(_1307_));
 NAND2_X1 _4332_ (.A1(_1307_),
    .A2(_1617_),
    .ZN(_1308_));
 OAI21_X1 _4333_ (.A(_1308_),
    .B1(_1617_),
    .B2(_1284_),
    .ZN(_1309_));
 MUX2_X1 _4334_ (.A(_1309_),
    .B(_1289_),
    .S(net88),
    .Z(_1310_));
 NOR2_X2 _4335_ (.A1(net140),
    .A2(_1264_),
    .ZN(_1311_));
 OAI21_X1 _4336_ (.A(_1306_),
    .B1(_1275_),
    .B2(_1311_),
    .ZN(_1312_));
 NAND2_X1 _4337_ (.A1(_1298_),
    .A2(_1312_),
    .ZN(_1313_));
 INV_X1 _4338_ (.A(_1313_),
    .ZN(_1314_));
 NAND3_X1 _4339_ (.A1(_1764_),
    .A2(net95),
    .A3(net128),
    .ZN(_1315_));
 NAND3_X1 _4340_ (.A1(_1755_),
    .A2(_1617_),
    .A3(net128),
    .ZN(_1316_));
 NAND3_X1 _4341_ (.A1(_1315_),
    .A2(_1303_),
    .A3(_1316_),
    .ZN(_1317_));
 AOI21_X1 _4342_ (.A(_1317_),
    .B1(_1250_),
    .B2(_2363_),
    .ZN(_1318_));
 AND2_X1 _4343_ (.A1(_1271_),
    .A2(_1273_),
    .ZN(_1319_));
 NAND2_X1 _4344_ (.A1(_1292_),
    .A2(_1293_),
    .ZN(_1320_));
 OAI21_X1 _4345_ (.A(_1252_),
    .B1(_1319_),
    .B2(_1320_),
    .ZN(_1321_));
 NAND2_X1 _4346_ (.A1(_1318_),
    .A2(_1321_),
    .ZN(_1322_));
 INV_X1 _4347_ (.A(_1322_),
    .ZN(_1323_));
 NAND3_X1 _4348_ (.A1(_1265_),
    .A2(_1314_),
    .A3(_1323_),
    .ZN(_1324_));
 NAND2_X1 _4349_ (.A1(_1244_),
    .A2(_1857_),
    .ZN(_1325_));
 NAND2_X1 _4350_ (.A1(_1325_),
    .A2(_1617_),
    .ZN(_1326_));
 NAND2_X1 _4351_ (.A1(_1244_),
    .A2(_1855_),
    .ZN(_1327_));
 INV_X1 _4352_ (.A(_1327_),
    .ZN(_1328_));
 OAI21_X1 _4353_ (.A(_1326_),
    .B1(_1328_),
    .B2(_1617_),
    .ZN(_1329_));
 OR2_X1 _4354_ (.A1(_1329_),
    .A2(_1252_),
    .ZN(_1330_));
 NAND2_X1 _4355_ (.A1(net134),
    .A2(_1871_),
    .ZN(_1331_));
 NAND2_X1 _4356_ (.A1(_1331_),
    .A2(net91),
    .ZN(_1332_));
 NOR2_X1 _4357_ (.A1(net135),
    .A2(_1876_),
    .ZN(_1333_));
 OAI21_X2 _4358_ (.A(_1332_),
    .B1(_1333_),
    .B2(net91),
    .ZN(_1334_));
 OAI21_X1 _4359_ (.A(_1330_),
    .B1(net88),
    .B2(_1334_),
    .ZN(_1335_));
 NAND2_X1 _4360_ (.A1(_1333_),
    .A2(net91),
    .ZN(_1336_));
 NAND2_X1 _4361_ (.A1(_1244_),
    .A2(_1901_),
    .ZN(_1337_));
 OAI21_X1 _4362_ (.A(_1336_),
    .B1(net91),
    .B2(_1337_),
    .ZN(_1338_));
 NAND2_X1 _4363_ (.A1(_1338_),
    .A2(net88),
    .ZN(_1339_));
 NAND2_X1 _4364_ (.A1(_1244_),
    .A2(_1905_),
    .ZN(_1340_));
 NAND2_X1 _4365_ (.A1(_1340_),
    .A2(net91),
    .ZN(_1341_));
 NOR2_X1 _4366_ (.A1(net135),
    .A2(_1920_),
    .ZN(_1342_));
 OAI21_X1 _4367_ (.A(_1341_),
    .B1(net91),
    .B2(_1342_),
    .ZN(_1343_));
 OAI21_X1 _4368_ (.A(_1339_),
    .B1(net88),
    .B2(_1343_),
    .ZN(_1344_));
 NOR2_X1 _4369_ (.A1(_1335_),
    .A2(_1344_),
    .ZN(_1345_));
 NOR2_X1 _4370_ (.A1(_1345_),
    .A2(_1264_),
    .ZN(_1346_));
 MUX2_X1 _4371_ (.A(_1340_),
    .B(_1337_),
    .S(net91),
    .Z(_1347_));
 INV_X1 _4372_ (.A(_1338_),
    .ZN(_1348_));
 NAND3_X1 _4373_ (.A1(_1347_),
    .A2(_1252_),
    .A3(_1348_),
    .ZN(_1349_));
 NAND2_X1 _4374_ (.A1(_1331_),
    .A2(_1617_),
    .ZN(_1350_));
 NAND2_X1 _4375_ (.A1(_1325_),
    .A2(net92),
    .ZN(_1351_));
 NAND2_X1 _4376_ (.A1(_1350_),
    .A2(_1351_),
    .ZN(_1352_));
 NAND3_X2 _4377_ (.A1(_1334_),
    .A2(net88),
    .A3(_1352_),
    .ZN(_1353_));
 NAND3_X2 _4378_ (.A1(_1349_),
    .A2(_1353_),
    .A3(_1264_),
    .ZN(_1354_));
 OAI21_X1 _4379_ (.A(_1617_),
    .B1(net135),
    .B2(_1923_),
    .ZN(_1355_));
 OAI21_X1 _4380_ (.A(_1355_),
    .B1(_1617_),
    .B2(_1342_),
    .ZN(_1356_));
 NAND3_X1 _4381_ (.A1(_1343_),
    .A2(_1356_),
    .A3(net88),
    .ZN(_1357_));
 NOR2_X1 _4382_ (.A1(net122),
    .A2(_1923_),
    .ZN(_1358_));
 NAND2_X1 _4383_ (.A1(_1358_),
    .A2(net91),
    .ZN(_1359_));
 OAI21_X2 _4384_ (.A(_1359_),
    .B1(net91),
    .B2(_1299_),
    .ZN(_1360_));
 OAI21_X1 _4385_ (.A(_1252_),
    .B1(_1299_),
    .B2(_1617_),
    .ZN(_1361_));
 OAI21_X2 _4386_ (.A(_1357_),
    .B1(_1360_),
    .B2(_1361_),
    .ZN(_1362_));
 OAI21_X2 _4387_ (.A(_1354_),
    .B1(_1362_),
    .B2(_1264_),
    .ZN(_1363_));
 NAND2_X1 _4388_ (.A1(_1307_),
    .A2(net93),
    .ZN(_1364_));
 OAI21_X1 _4389_ (.A(_1364_),
    .B1(net93),
    .B2(_1328_),
    .ZN(_1365_));
 MUX2_X1 _4390_ (.A(_1352_),
    .B(_1365_),
    .S(net88),
    .Z(_1366_));
 AOI21_X1 _4391_ (.A(net141),
    .B1(_1310_),
    .B2(_1366_),
    .ZN(_1367_));
 NOR3_X2 _4392_ (.A1(_1346_),
    .A2(_1363_),
    .A3(_1367_),
    .ZN(_1368_));
 NOR2_X1 _4393_ (.A1(_1362_),
    .A2(net144),
    .ZN(_1369_));
 NAND2_X1 _4394_ (.A1(net88),
    .A2(_1360_),
    .ZN(_1370_));
 NOR2_X2 _4395_ (.A1(_1370_),
    .A2(net144),
    .ZN(_1371_));
 NOR4_X1 _4396_ (.A1(_1369_),
    .A2(_1371_),
    .A3(_1303_),
    .A4(_1301_),
    .ZN(_1372_));
 NOR2_X1 _4397_ (.A1(_1286_),
    .A2(net141),
    .ZN(_1373_));
 NAND3_X1 _4398_ (.A1(_1285_),
    .A2(_1309_),
    .A3(net88),
    .ZN(_1374_));
 NAND3_X1 _4399_ (.A1(_1329_),
    .A2(_1365_),
    .A3(_1252_),
    .ZN(_1375_));
 NAND2_X1 _4400_ (.A1(_1374_),
    .A2(_1375_),
    .ZN(_1376_));
 NAND2_X1 _4401_ (.A1(_1373_),
    .A2(_1376_),
    .ZN(_1377_));
 NAND2_X1 _4402_ (.A1(_1349_),
    .A2(_1353_),
    .ZN(_1378_));
 NAND3_X1 _4403_ (.A1(_1366_),
    .A2(_1378_),
    .A3(net142),
    .ZN(_1379_));
 NAND2_X1 _4404_ (.A1(_1377_),
    .A2(_1379_),
    .ZN(_1380_));
 NAND2_X2 _4405_ (.A1(net133),
    .A2(net88),
    .ZN(_1381_));
 INV_X1 _4406_ (.A(_1356_),
    .ZN(_1382_));
 OAI21_X2 _4407_ (.A(_1381_),
    .B1(_1382_),
    .B2(net88),
    .ZN(_1383_));
 NAND2_X1 _4408_ (.A1(_1383_),
    .A2(net143),
    .ZN(_1384_));
 OAI21_X1 _4409_ (.A(_1384_),
    .B1(_1335_),
    .B2(net143),
    .ZN(_1385_));
 INV_X1 _4410_ (.A(_1385_),
    .ZN(_1386_));
 NAND2_X1 _4411_ (.A1(_1386_),
    .A2(_1306_),
    .ZN(_1387_));
 NAND4_X1 _4412_ (.A1(_1368_),
    .A2(_1372_),
    .A3(_1380_),
    .A4(_1387_),
    .ZN(_1388_));
 NAND2_X1 _4413_ (.A1(_1324_),
    .A2(_1388_),
    .ZN(_1389_));
 NAND3_X1 _4414_ (.A1(_1368_),
    .A2(_1380_),
    .A3(_1385_),
    .ZN(_1390_));
 NAND2_X1 _4415_ (.A1(_1390_),
    .A2(_1303_),
    .ZN(_1391_));
 OR2_X1 _4416_ (.A1(_1295_),
    .A2(_2372_),
    .ZN(_1392_));
 NAND2_X1 _4417_ (.A1(_1383_),
    .A2(_1264_),
    .ZN(_1393_));
 OAI21_X1 _4418_ (.A(_1393_),
    .B1(_1264_),
    .B2(_1300_),
    .ZN(_1394_));
 NAND2_X1 _4419_ (.A1(_1370_),
    .A2(net143),
    .ZN(_1395_));
 OAI21_X1 _4420_ (.A(_1395_),
    .B1(_1344_),
    .B2(net143),
    .ZN(_1396_));
 NAND2_X1 _4421_ (.A1(_1396_),
    .A2(_1394_),
    .ZN(_1397_));
 INV_X1 _4422_ (.A(_1397_),
    .ZN(_1398_));
 NAND2_X1 _4423_ (.A1(_1371_),
    .A2(_1303_),
    .ZN(_1399_));
 NAND3_X1 _4424_ (.A1(_1399_),
    .A2(_2376_),
    .A3(_1304_),
    .ZN(_1400_));
 NOR2_X1 _4425_ (.A1(_1376_),
    .A2(_1264_),
    .ZN(_1401_));
 NOR2_X1 _4426_ (.A1(_1400_),
    .A2(_1401_),
    .ZN(_1402_));
 NAND2_X1 _4427_ (.A1(_1369_),
    .A2(_1303_),
    .ZN(_1403_));
 NAND4_X1 _4428_ (.A1(_1392_),
    .A2(_1398_),
    .A3(_1402_),
    .A4(_1403_),
    .ZN(_1404_));
 INV_X1 _4429_ (.A(_1404_),
    .ZN(_1405_));
 NAND2_X1 _4430_ (.A1(_1391_),
    .A2(_1405_),
    .ZN(_1406_));
 INV_X1 _4431_ (.A(_1406_),
    .ZN(_1407_));
 NAND2_X1 _4432_ (.A1(_1389_),
    .A2(_1407_),
    .ZN(_1408_));
 XOR2_X1 _4433_ (.A(net138),
    .B(_2375_),
    .Z(_1409_));
 OAI21_X1 _4434_ (.A(_1303_),
    .B1(_1397_),
    .B2(_1363_),
    .ZN(_1410_));
 NAND4_X1 _4435_ (.A1(_1403_),
    .A2(_1305_),
    .A3(_1304_),
    .A4(_1399_),
    .ZN(_1411_));
 INV_X1 _4436_ (.A(_1411_),
    .ZN(_1412_));
 AOI21_X1 _4437_ (.A(_1409_),
    .B1(_1410_),
    .B2(_1412_),
    .ZN(_1413_));
 NAND2_X2 _4438_ (.A1(_1408_),
    .A2(_1413_),
    .ZN(_1414_));
 INV_X1 _4439_ (.A(_2356_),
    .ZN(_1415_));
 NAND3_X1 _4440_ (.A1(_1643_),
    .A2(_2364_),
    .A3(_1553_),
    .ZN(_1416_));
 OAI21_X1 _4441_ (.A(_1571_),
    .B1(_1884_),
    .B2(_1416_),
    .ZN(_1417_));
 NOR2_X1 _4442_ (.A1(_1415_),
    .A2(_1417_),
    .ZN(_1418_));
 NAND2_X2 _4443_ (.A1(_1414_),
    .A2(_1418_),
    .ZN(_1419_));
 OR4_X1 _4444_ (.A1(_1755_),
    .A2(_1778_),
    .A3(_1769_),
    .A4(_1764_),
    .ZN(_1420_));
 NOR4_X1 _4445_ (.A1(_1291_),
    .A2(_1749_),
    .A3(_1742_),
    .A4(_1824_),
    .ZN(_1421_));
 NOR4_X1 _4446_ (.A1(_1905_),
    .A2(_1924_),
    .A3(_1919_),
    .A4(_1200_),
    .ZN(_1422_));
 NOR4_X1 _4447_ (.A1(_1857_),
    .A2(_1875_),
    .A3(_1871_),
    .A4(_1901_),
    .ZN(_1423_));
 NOR4_X1 _4448_ (.A1(_1820_),
    .A2(_1816_),
    .A3(_1827_),
    .A4(_1855_),
    .ZN(_1424_));
 NAND4_X1 _4449_ (.A1(_1421_),
    .A2(_1422_),
    .A3(_1423_),
    .A4(_1424_),
    .ZN(_1425_));
 NAND4_X1 _4450_ (.A1(_1781_),
    .A2(_1798_),
    .A3(_1259_),
    .A4(_1633_),
    .ZN(_1426_));
 OR4_X1 _4451_ (.A1(_1418_),
    .A2(_1420_),
    .A3(_1425_),
    .A4(_1426_),
    .ZN(_1427_));
 NAND2_X1 _4452_ (.A1(_1419_),
    .A2(_1427_),
    .ZN(_1428_));
 NAND2_X1 _4453_ (.A1(_1428_),
    .A2(_1627_),
    .ZN(_1429_));
 NAND3_X1 _4454_ (.A1(_1419_),
    .A2(_1733_),
    .A3(_1427_),
    .ZN(_1430_));
 NAND2_X1 _4455_ (.A1(_1430_),
    .A2(_1429_),
    .ZN(_1431_));
 INV_X1 _4456_ (.A(_1431_),
    .ZN(_2039_));
 INV_X1 _4457_ (.A(_0064_),
    .ZN(_1981_));
 INV_X1 _4458_ (.A(_2059_),
    .ZN(_2100_));
 INV_X1 _4459_ (.A(_1090_),
    .ZN(_2043_));
 NOR2_X1 _4460_ (.A1(net150),
    .A2(_0242_),
    .ZN(_2122_));
 NOR2_X4 _4461_ (.A1(_0991_),
    .A2(_1081_),
    .ZN(_2044_));
 INV_X1 _4462_ (.A(_2091_),
    .ZN(_2052_));
 INV_X1 _4463_ (.A(_2140_),
    .ZN(_1432_));
 INV_X1 _4464_ (.A(_2141_),
    .ZN(_1433_));
 INV_X1 _4465_ (.A(_2137_),
    .ZN(_1434_));
 NAND2_X1 _4466_ (.A1(_2138_),
    .A2(_2141_),
    .ZN(_1435_));
 OAI221_X2 _4467_ (.A(_1432_),
    .B1(_1433_),
    .B2(_1434_),
    .C1(_2056_),
    .C2(_1435_),
    .ZN(_2061_));
 INV_X1 _4468_ (.A(_1067_),
    .ZN(_2180_));
 INV_X1 _4469_ (.A(_2184_),
    .ZN(_1436_));
 INV_X1 _4470_ (.A(_1080_),
    .ZN(_1437_));
 NOR2_X2 _4471_ (.A1(_1436_),
    .A2(_1437_),
    .ZN(_2188_));
 INV_X1 _4472_ (.A(_1946_),
    .ZN(_1950_));
 INV_X1 _4473_ (.A(_2227_),
    .ZN(_2231_));
 NAND2_X1 _4474_ (.A1(_1176_),
    .A2(_1565_),
    .ZN(_1438_));
 XNOR2_X1 _4475_ (.A(_1733_),
    .B(_1438_),
    .ZN(_2273_));
 NAND2_X1 _4476_ (.A1(_1885_),
    .A2(_1565_),
    .ZN(_1439_));
 XNOR2_X1 _4477_ (.A(_1627_),
    .B(_1439_),
    .ZN(_1440_));
 INV_X1 _4478_ (.A(_1440_),
    .ZN(_1978_));
 NOR2_X1 _4479_ (.A1(_1134_),
    .A2(_1643_),
    .ZN(_1441_));
 NAND2_X1 _4480_ (.A1(_1441_),
    .A2(_1565_),
    .ZN(_1442_));
 XNOR2_X1 _4481_ (.A(_1733_),
    .B(_1442_),
    .ZN(_2279_));
 NAND2_X1 _4482_ (.A1(_1892_),
    .A2(_1565_),
    .ZN(_1443_));
 XNOR2_X1 _4483_ (.A(_1627_),
    .B(_1443_),
    .ZN(_1444_));
 INV_X1 _4484_ (.A(_1444_),
    .ZN(_1983_));
 NOR2_X1 _4485_ (.A1(net90),
    .A2(net26),
    .ZN(_1445_));
 AOI21_X1 _4486_ (.A(_1445_),
    .B1(_2252_),
    .B2(net90),
    .ZN(_1446_));
 XNOR2_X1 _4487_ (.A(_1648_),
    .B(_1446_),
    .ZN(_2285_));
 NOR2_X1 _4488_ (.A1(net90),
    .A2(net25),
    .ZN(_1447_));
 AOI21_X1 _4489_ (.A(_1447_),
    .B1(_2255_),
    .B2(net90),
    .ZN(_1448_));
 XNOR2_X2 _4490_ (.A(_1648_),
    .B(_1448_),
    .ZN(_1988_));
 NOR2_X1 _4491_ (.A1(_1216_),
    .A2(_1814_),
    .ZN(_1449_));
 XNOR2_X1 _4492_ (.A(_1733_),
    .B(_1449_),
    .ZN(_1450_));
 INV_X1 _4493_ (.A(_1450_),
    .ZN(_2291_));
 NAND2_X1 _4494_ (.A1(_1221_),
    .A2(_1565_),
    .ZN(_1451_));
 XNOR2_X1 _4495_ (.A(_1451_),
    .B(_1627_),
    .ZN(_1452_));
 INV_X1 _4496_ (.A(_1452_),
    .ZN(_1993_));
 NAND3_X1 _4497_ (.A1(_1231_),
    .A2(_1565_),
    .A3(_1232_),
    .ZN(_1453_));
 XNOR2_X1 _4498_ (.A(_1627_),
    .B(_1453_),
    .ZN(_1454_));
 INV_X1 _4499_ (.A(_1454_),
    .ZN(_2297_));
 INV_X1 _4500_ (.A(_1998_),
    .ZN(_2301_));
 NOR2_X1 _4501_ (.A1(net90),
    .A2(_1823_),
    .ZN(_1455_));
 XNOR2_X1 _4502_ (.A(_1648_),
    .B(_1455_),
    .ZN(_2305_));
 AOI21_X1 _4503_ (.A(_1814_),
    .B1(_1895_),
    .B2(net89),
    .ZN(_1456_));
 NAND2_X1 _4504_ (.A1(_1891_),
    .A2(_1643_),
    .ZN(_1457_));
 NAND2_X1 _4505_ (.A1(_1456_),
    .A2(_1457_),
    .ZN(_1458_));
 XNOR2_X1 _4506_ (.A(_1458_),
    .B(_1627_),
    .ZN(_1459_));
 INV_X1 _4507_ (.A(_1459_),
    .ZN(_2003_));
 NAND2_X1 _4508_ (.A1(_1121_),
    .A2(_1643_),
    .ZN(_1460_));
 NAND2_X1 _4509_ (.A1(_1180_),
    .A2(net89),
    .ZN(_1461_));
 NAND3_X1 _4510_ (.A1(_1460_),
    .A2(_1461_),
    .A3(_1565_),
    .ZN(_1462_));
 XNOR2_X1 _4511_ (.A(_1462_),
    .B(_1627_),
    .ZN(_1463_));
 INV_X1 _4512_ (.A(_1463_),
    .ZN(_2311_));
 INV_X1 _4513_ (.A(_2008_),
    .ZN(_2315_));
 AOI21_X1 _4514_ (.A(net89),
    .B1(_1213_),
    .B2(_1215_),
    .ZN(_1464_));
 OAI21_X1 _4515_ (.A(_1565_),
    .B1(_1211_),
    .B2(_1643_),
    .ZN(_1465_));
 NOR2_X1 _4516_ (.A1(_1464_),
    .A2(_1465_),
    .ZN(_1466_));
 XNOR2_X1 _4517_ (.A(_1733_),
    .B(_1466_),
    .ZN(_1467_));
 INV_X1 _4518_ (.A(_1467_),
    .ZN(_2319_));
 INV_X1 _4519_ (.A(_2013_),
    .ZN(_2323_));
 NOR2_X1 _4520_ (.A1(net90),
    .A2(_1870_),
    .ZN(_1468_));
 XNOR2_X1 _4521_ (.A(_1648_),
    .B(_1468_),
    .ZN(_2327_));
 INV_X1 _4522_ (.A(_2018_),
    .ZN(_2331_));
 NAND2_X1 _4523_ (.A1(_1441_),
    .A2(_1843_),
    .ZN(_1469_));
 NAND3_X1 _4524_ (.A1(_1140_),
    .A2(_1643_),
    .A3(_1148_),
    .ZN(_1470_));
 NAND2_X1 _4525_ (.A1(_1208_),
    .A2(_1576_),
    .ZN(_1471_));
 OAI21_X1 _4526_ (.A(_1471_),
    .B1(_1198_),
    .B2(_1576_),
    .ZN(_1472_));
 AOI21_X1 _4527_ (.A(_1814_),
    .B1(_1472_),
    .B2(net89),
    .ZN(_1473_));
 NAND2_X1 _4528_ (.A1(_1470_),
    .A2(_1473_),
    .ZN(_1474_));
 NAND2_X1 _4529_ (.A1(_1469_),
    .A2(_1474_),
    .ZN(_1475_));
 XNOR2_X1 _4530_ (.A(_1733_),
    .B(_1475_),
    .ZN(_1476_));
 INV_X1 _4531_ (.A(_1476_),
    .ZN(_2335_));
 INV_X1 _4532_ (.A(_2022_),
    .ZN(_2339_));
 NOR2_X1 _4533_ (.A1(net90),
    .A2(_1918_),
    .ZN(_1477_));
 XNOR2_X1 _4534_ (.A(_1648_),
    .B(_1477_),
    .ZN(_2343_));
 INV_X1 _4535_ (.A(_2027_),
    .ZN(_2347_));
 NOR2_X1 _4536_ (.A1(net90),
    .A2(_1199_),
    .ZN(_1478_));
 XNOR2_X1 _4537_ (.A(_1648_),
    .B(_1478_),
    .ZN(_2351_));
 FA_X1 _4538_ (.A(net33),
    .B(_1937_),
    .CI(_1938_),
    .CO(_1939_),
    .S(_1940_));
 FA_X1 _4539_ (.A(_1941_),
    .B(_1942_),
    .CI(_1943_),
    .CO(_1944_),
    .S(_1945_));
 FA_X1 _4540_ (.A(net34),
    .B(_1946_),
    .CI(_1939_),
    .CO(_1947_),
    .S(_1948_));
 FA_X1 _4541_ (.A(_1949_),
    .B(_1950_),
    .CI(_1944_),
    .CO(_1951_),
    .S(_1952_));
 FA_X1 _4542_ (.A(_1953_),
    .B(_1954_),
    .CI(_1955_),
    .CO(_1956_),
    .S(_1957_));
 FA_X1 _4543_ (.A(net36),
    .B(_1958_),
    .CI(_1959_),
    .CO(_1960_),
    .S(_1961_));
 FA_X1 _4544_ (.A(net38),
    .B(_1962_),
    .CI(_1963_),
    .CO(_1964_),
    .S(_1965_));
 FA_X1 _4545_ (.A(_1966_),
    .B(_1967_),
    .CI(_1968_),
    .CO(_1969_),
    .S(_1970_));
 FA_X1 _4546_ (.A(_1971_),
    .B(_1972_),
    .CI(_1973_),
    .CO(_1974_),
    .S(_1975_));
 FA_X1 _4547_ (.A(net146),
    .B(_1977_),
    .CI(_1978_),
    .CO(_1979_),
    .S(_1980_));
 FA_X1 _4548_ (.A(_1981_),
    .B(_1982_),
    .CI(_1983_),
    .CO(_1984_),
    .S(_1985_));
 FA_X1 _4549_ (.A(_1986_),
    .B(_1987_),
    .CI(_1988_),
    .CO(_1989_),
    .S(_1990_));
 FA_X1 _4550_ (.A(_1991_),
    .B(_1992_),
    .CI(_1993_),
    .CO(_1994_),
    .S(_1995_));
 FA_X1 _4551_ (.A(_1996_),
    .B(_1997_),
    .CI(_1998_),
    .CO(_1999_),
    .S(_2000_));
 FA_X1 _4552_ (.A(_2001_),
    .B(_2002_),
    .CI(_2003_),
    .CO(_2004_),
    .S(_2005_));
 FA_X1 _4553_ (.A(_2006_),
    .B(_2007_),
    .CI(_2008_),
    .CO(_2009_),
    .S(_2010_));
 FA_X1 _4554_ (.A(_2011_),
    .B(_2012_),
    .CI(_2013_),
    .CO(_2014_),
    .S(_2015_));
 FA_X1 _4555_ (.A(net130),
    .B(_2017_),
    .CI(_2018_),
    .CO(_2019_),
    .S(_2020_));
 FA_X1 _4556_ (.A(_2021_),
    .B(_2022_),
    .CI(_2023_),
    .CO(_2024_),
    .S(_2025_));
 FA_X1 _4557_ (.A(_2026_),
    .B(_2027_),
    .CI(net119),
    .CO(_2029_),
    .S(_2030_));
 FA_X1 _4558_ (.A(_2031_),
    .B(_2032_),
    .CI(_2033_),
    .CO(_2034_),
    .S(_2035_));
 FA_X1 _4559_ (.A(_2036_),
    .B(_2037_),
    .CI(_2033_),
    .CO(_2031_),
    .S(_2038_));
 FA_X1 _4560_ (.A(_2039_),
    .B(_2033_),
    .CI(_2040_),
    .CO(_2036_),
    .S(_2041_));
 FA_X1 _4561_ (.A(_2042_),
    .B(_2043_),
    .CI(_2044_),
    .CO(_2045_),
    .S(_2046_));
 FA_X1 _4562_ (.A(_2047_),
    .B(_2048_),
    .CI(_2045_),
    .CO(_2049_),
    .S(_2050_));
 FA_X1 _4563_ (.A(net107),
    .B(_2052_),
    .CI(_2049_),
    .CO(_2053_),
    .S(_2054_));
 FA_X1 _4564_ (.A(_2055_),
    .B(_2056_),
    .CI(_2057_),
    .CO(_2058_),
    .S(net68));
 FA_X1 _4565_ (.A(_2059_),
    .B(_2060_),
    .CI(_2061_),
    .CO(_2062_),
    .S(_2063_));
 HA_X1 _4566_ (.A(_2064_),
    .B(_2065_),
    .CO(_2066_),
    .S(_2067_));
 HA_X1 _4567_ (.A(_2068_),
    .B(_2069_),
    .CO(_2070_),
    .S(_2071_));
 HA_X1 _4568_ (.A(_2072_),
    .B(_2073_),
    .CO(_2074_),
    .S(_2075_));
 HA_X1 _4569_ (.A(_2076_),
    .B(_2077_),
    .CO(_2078_),
    .S(_2079_));
 HA_X1 _4570_ (.A(_2080_),
    .B(_2081_),
    .CO(_2082_),
    .S(_2051_));
 HA_X1 _4571_ (.A(_2083_),
    .B(_2084_),
    .CO(_2085_),
    .S(_2086_));
 HA_X1 _4572_ (.A(_2087_),
    .B(_2088_),
    .CO(_2089_),
    .S(_2090_));
 HA_X1 _4573_ (.A(_2087_),
    .B(_2088_),
    .CO(_2091_),
    .S(_2092_));
 HA_X1 _4574_ (.A(_2043_),
    .B(_2093_),
    .CO(_2094_),
    .S(_2095_));
 HA_X1 _4575_ (.A(_2096_),
    .B(_2081_),
    .CO(_2097_),
    .S(_2098_));
 HA_X1 _4576_ (.A(_2099_),
    .B(_2100_),
    .CO(_2101_),
    .S(_2102_));
 HA_X1 _4577_ (.A(_2103_),
    .B(_2065_),
    .CO(_2104_),
    .S(_2105_));
 HA_X1 _4578_ (.A(_2106_),
    .B(_2043_),
    .CO(_2107_),
    .S(_2108_));
 HA_X1 _4579_ (.A(_2107_),
    .B(_2109_),
    .CO(_2096_),
    .S(_2110_));
 HA_X1 _4580_ (.A(_2111_),
    .B(_0295_),
    .CO(_2113_),
    .S(_2114_));
 HA_X1 _4581_ (.A(_2111_),
    .B(_0232_),
    .CO(_2116_),
    .S(_2117_));
 HA_X1 _4582_ (.A(_2116_),
    .B(_2118_),
    .CO(_2119_),
    .S(_2120_));
 HA_X1 _4583_ (.A(_2121_),
    .B(_2122_),
    .CO(_2123_),
    .S(_2124_));
 HA_X1 _4584_ (.A(_2125_),
    .B(_2126_),
    .CO(_2127_),
    .S(_2128_));
 HA_X1 _4585_ (.A(_2129_),
    .B(_2130_),
    .CO(_2131_),
    .S(_2132_));
 HA_X1 _4586_ (.A(_2093_),
    .B(_2046_),
    .CO(_2048_),
    .S(net64));
 HA_X1 _4587_ (.A(net106),
    .B(_2052_),
    .CO(_2133_),
    .S(_2134_));
 HA_X1 _4588_ (.A(_2075_),
    .B(_2082_),
    .CO(_2135_),
    .S(_2136_));
 HA_X1 _4589_ (.A(_2067_),
    .B(_2074_),
    .CO(_2137_),
    .S(_2138_));
 HA_X1 _4590_ (.A(_2139_),
    .B(_2066_),
    .CO(_2140_),
    .S(_2141_));
 HA_X1 _4591_ (.A(_2142_),
    .B(_2059_),
    .CO(_2143_),
    .S(_2144_));
 HA_X1 _4592_ (.A(_2145_),
    .B(_2100_),
    .CO(_2146_),
    .S(_2147_));
 HA_X1 _4593_ (.A(_2148_),
    .B(_2149_),
    .CO(_2150_),
    .S(_2151_));
 HA_X1 _4594_ (.A(_2150_),
    .B(_2152_),
    .CO(_2153_),
    .S(_2154_));
 HA_X1 _4595_ (.A(_2155_),
    .B(_2156_),
    .CO(_2157_),
    .S(_2158_));
 HA_X1 _4596_ (.A(_2159_),
    .B(_2160_),
    .CO(_2161_),
    .S(_2162_));
 HA_X1 _4597_ (.A(_2163_),
    .B(_2164_),
    .CO(_2165_),
    .S(_2166_));
 HA_X1 _4598_ (.A(_2167_),
    .B(_2168_),
    .CO(_2169_),
    .S(_2170_));
 HA_X1 _4599_ (.A(_2171_),
    .B(_2172_),
    .CO(_2173_),
    .S(_2174_));
 HA_X1 _4600_ (.A(_2175_),
    .B(_2176_),
    .CO(_2177_),
    .S(_2178_));
 HA_X1 _4601_ (.A(_2179_),
    .B(_2180_),
    .CO(_2181_),
    .S(_2182_));
 HA_X1 _4602_ (.A(_2183_),
    .B(_2184_),
    .CO(_2185_),
    .S(_2186_));
 HA_X1 _4603_ (.A(_2187_),
    .B(_2188_),
    .CO(_2189_),
    .S(_2190_));
 HA_X1 _4604_ (.A(_2191_),
    .B(_2192_),
    .CO(_2193_),
    .S(_2194_));
 HA_X1 _4605_ (.A(_2195_),
    .B(net40),
    .CO(_2196_),
    .S(_2197_));
 HA_X1 _4606_ (.A(_1966_),
    .B(_1967_),
    .CO(_2198_),
    .S(_2199_));
 HA_X1 _4607_ (.A(net38),
    .B(_1962_),
    .CO(_2200_),
    .S(_2201_));
 HA_X1 _4608_ (.A(_2202_),
    .B(_1967_),
    .CO(_2203_),
    .S(_2204_));
 HA_X1 _4609_ (.A(net37),
    .B(_1962_),
    .CO(_2205_),
    .S(_2206_));
 HA_X1 _4610_ (.A(_1953_),
    .B(_1954_),
    .CO(_2207_),
    .S(_2208_));
 HA_X1 _4611_ (.A(net36),
    .B(_1958_),
    .CO(_2209_),
    .S(_2210_));
 HA_X1 _4612_ (.A(_2211_),
    .B(_2212_),
    .CO(_2213_),
    .S(_2214_));
 HA_X1 _4613_ (.A(net35),
    .B(_2215_),
    .CO(_2216_),
    .S(_2217_));
 HA_X1 _4614_ (.A(_2218_),
    .B(_2219_),
    .CO(_2220_),
    .S(_2221_));
 HA_X1 _4615_ (.A(_1949_),
    .B(_1950_),
    .CO(_2222_),
    .S(_2223_));
 HA_X1 _4616_ (.A(net34),
    .B(_1946_),
    .CO(_2224_),
    .S(_2225_));
 HA_X1 _4617_ (.A(_2226_),
    .B(_2227_),
    .CO(_2228_),
    .S(_2229_));
 HA_X1 _4618_ (.A(_1505_),
    .B(_2231_),
    .CO(_2218_),
    .S(_2232_));
 HA_X1 _4619_ (.A(_2233_),
    .B(_2234_),
    .CO(_2235_),
    .S(_2236_));
 HA_X1 _4620_ (.A(_2237_),
    .B(_2228_),
    .CO(_2238_),
    .S(_2239_));
 HA_X1 _4621_ (.A(net31),
    .B(_2240_),
    .CO(_2241_),
    .S(_2242_));
 HA_X1 _4622_ (.A(net30),
    .B(_2243_),
    .CO(_2244_),
    .S(_2245_));
 HA_X1 _4623_ (.A(net29),
    .B(_2246_),
    .CO(_2247_),
    .S(_2248_));
 HA_X1 _4624_ (.A(net27),
    .B(_2249_),
    .CO(_2250_),
    .S(_2251_));
 HA_X1 _4625_ (.A(net26),
    .B(_2252_),
    .CO(_2253_),
    .S(_2254_));
 HA_X1 _4626_ (.A(net25),
    .B(_2255_),
    .CO(_2256_),
    .S(_2257_));
 HA_X1 _4627_ (.A(net24),
    .B(_2258_),
    .CO(_2259_),
    .S(_2260_));
 HA_X1 _4628_ (.A(net23),
    .B(_2261_),
    .CO(_2262_),
    .S(_2263_));
 HA_X1 _4629_ (.A(net22),
    .B(_2264_),
    .CO(_2265_),
    .S(_2266_));
 HA_X1 _4630_ (.A(_2267_),
    .B(_2268_),
    .CO(_1943_),
    .S(_2269_));
 HA_X1 _4631_ (.A(net32),
    .B(_2270_),
    .CO(_1937_),
    .S(_2271_));
 HA_X1 _4632_ (.A(_2272_),
    .B(_2273_),
    .CO(_2274_),
    .S(_2275_));
 HA_X1 _4633_ (.A(_1977_),
    .B(_1978_),
    .CO(_2276_),
    .S(_2277_));
 HA_X1 _4634_ (.A(_2278_),
    .B(_2279_),
    .CO(_2280_),
    .S(_2281_));
 HA_X1 _4635_ (.A(_1982_),
    .B(_1983_),
    .CO(_2282_),
    .S(_2283_));
 HA_X1 _4636_ (.A(_2284_),
    .B(_2285_),
    .CO(_2286_),
    .S(_2287_));
 HA_X1 _4637_ (.A(_1987_),
    .B(_1988_),
    .CO(_2288_),
    .S(_2289_));
 HA_X1 _4638_ (.A(_2290_),
    .B(_2291_),
    .CO(_2292_),
    .S(_2293_));
 HA_X1 _4639_ (.A(_1992_),
    .B(_1993_),
    .CO(_2294_),
    .S(_2295_));
 HA_X1 _4640_ (.A(_2296_),
    .B(_2297_),
    .CO(_2298_),
    .S(_2299_));
 HA_X1 _4641_ (.A(_2300_),
    .B(_2301_),
    .CO(_2302_),
    .S(_2303_));
 HA_X1 _4642_ (.A(_2304_),
    .B(_2305_),
    .CO(_2306_),
    .S(_2307_));
 HA_X1 _4643_ (.A(_2002_),
    .B(_2003_),
    .CO(_2308_),
    .S(_2309_));
 HA_X1 _4644_ (.A(_2310_),
    .B(_2311_),
    .CO(_2312_),
    .S(_2313_));
 HA_X1 _4645_ (.A(_2314_),
    .B(_2315_),
    .CO(_2316_),
    .S(_2317_));
 HA_X1 _4646_ (.A(_2318_),
    .B(_2319_),
    .CO(_2320_),
    .S(_2321_));
 HA_X1 _4647_ (.A(_2322_),
    .B(_2323_),
    .CO(_2324_),
    .S(_2325_));
 HA_X1 _4648_ (.A(_2326_),
    .B(_2327_),
    .CO(_2328_),
    .S(_2329_));
 HA_X1 _4649_ (.A(_2330_),
    .B(_2331_),
    .CO(_2332_),
    .S(_2333_));
 HA_X1 _4650_ (.A(_2334_),
    .B(_2335_),
    .CO(_2336_),
    .S(_2337_));
 HA_X1 _4651_ (.A(_2338_),
    .B(_2339_),
    .CO(_2340_),
    .S(_2341_));
 HA_X1 _4652_ (.A(_2342_),
    .B(_2343_),
    .CO(_2344_),
    .S(_2345_));
 HA_X1 _4653_ (.A(_2346_),
    .B(_2347_),
    .CO(_2348_),
    .S(_2349_));
 HA_X1 _4654_ (.A(_2350_),
    .B(_2351_),
    .CO(_2352_),
    .S(_2353_));
 HA_X1 _4655_ (.A(_2032_),
    .B(_2033_),
    .CO(_2354_),
    .S(_2355_));
 HA_X1 _4656_ (.A(_2356_),
    .B(_2357_),
    .CO(_2358_),
    .S(_2359_));
 HA_X1 _4657_ (.A(_1617_),
    .B(_1620_),
    .CO(_2362_),
    .S(_2363_));
 HA_X1 _4658_ (.A(net94),
    .B(_1620_),
    .CO(_2364_),
    .S(_2365_));
 HA_X1 _4659_ (.A(_2269_),
    .B(_1546_),
    .CO(_2367_),
    .S(_2368_));
 HA_X1 _4660_ (.A(_1553_),
    .B(net139),
    .CO(_2371_),
    .S(_2372_));
 HA_X1 _4661_ (.A(net136),
    .B(_2374_),
    .CO(_2375_),
    .S(_2376_));
 TAPCELL_X1 PHY_0 ();
 BUF_X2 input11 (.A(operand_fp16_i[4]),
    .Z(net11));
 BUF_X2 input12 (.A(operand_fp16_i[5]),
    .Z(net12));
 BUF_X2 input13 (.A(operand_fp16_i[6]),
    .Z(net13));
 BUF_X4 input14 (.A(operand_fp16_i[7]),
    .Z(net14));
 BUF_X2 input15 (.A(operand_fp16_i[8]),
    .Z(net15));
 BUF_X2 input16 (.A(operand_fp16_i[9]),
    .Z(net16));
 BUF_X1 input17 (.A(operand_fp32_i[0]),
    .Z(net17));
 BUF_X1 input18 (.A(operand_fp32_i[10]),
    .Z(net18));
 BUF_X1 input19 (.A(operand_fp32_i[11]),
    .Z(net19));
 BUF_X1 input20 (.A(operand_fp32_i[12]),
    .Z(net20));
 BUF_X1 input21 (.A(operand_fp32_i[13]),
    .Z(net21));
 BUF_X1 input22 (.A(operand_fp32_i[14]),
    .Z(net22));
 BUF_X1 input23 (.A(operand_fp32_i[15]),
    .Z(net23));
 BUF_X1 input24 (.A(operand_fp32_i[16]),
    .Z(net24));
 BUF_X1 input25 (.A(operand_fp32_i[17]),
    .Z(net25));
 BUF_X1 input26 (.A(operand_fp32_i[18]),
    .Z(net26));
 BUF_X1 input27 (.A(operand_fp32_i[19]),
    .Z(net27));
 BUF_X1 input28 (.A(operand_fp32_i[1]),
    .Z(net28));
 BUF_X1 input29 (.A(operand_fp32_i[20]),
    .Z(net29));
 BUF_X1 input30 (.A(operand_fp32_i[21]),
    .Z(net30));
 BUF_X1 input31 (.A(operand_fp32_i[22]),
    .Z(net31));
 BUF_X1 input32 (.A(operand_fp32_i[23]),
    .Z(net32));
 BUF_X1 input33 (.A(operand_fp32_i[24]),
    .Z(net33));
 BUF_X2 input34 (.A(operand_fp32_i[25]),
    .Z(net34));
 BUF_X1 input35 (.A(operand_fp32_i[26]),
    .Z(net35));
 CLKBUF_X2 input36 (.A(operand_fp32_i[27]),
    .Z(net36));
 BUF_X1 input37 (.A(operand_fp32_i[28]),
    .Z(net37));
 BUF_X2 input38 (.A(operand_fp32_i[29]),
    .Z(net38));
 BUF_X1 input39 (.A(operand_fp32_i[2]),
    .Z(net39));
 BUF_X1 input40 (.A(operand_fp32_i[30]),
    .Z(net40));
 BUF_X1 input41 (.A(operand_fp32_i[31]),
    .Z(net41));
 BUF_X1 input42 (.A(operand_fp32_i[3]),
    .Z(net42));
 BUF_X1 input43 (.A(operand_fp32_i[4]),
    .Z(net43));
 BUF_X1 input44 (.A(operand_fp32_i[5]),
    .Z(net44));
 BUF_X1 input45 (.A(operand_fp32_i[6]),
    .Z(net45));
 BUF_X1 input46 (.A(operand_fp32_i[7]),
    .Z(net46));
 BUF_X1 input47 (.A(operand_fp32_i[8]),
    .Z(net47));
 BUF_X1 input48 (.A(operand_fp32_i[9]),
    .Z(net48));
 BUF_X1 output49 (.A(net49),
    .Z(result_o[0]));
 BUF_X1 output50 (.A(net50),
    .Z(result_o[10]));
 BUF_X1 output51 (.A(net51),
    .Z(result_o[11]));
 BUF_X1 output52 (.A(net52),
    .Z(result_o[12]));
 BUF_X1 output53 (.A(net53),
    .Z(result_o[13]));
 BUF_X1 output54 (.A(net54),
    .Z(result_o[14]));
 BUF_X1 output55 (.A(net55),
    .Z(result_o[15]));
 BUF_X1 output56 (.A(net56),
    .Z(result_o[16]));
 BUF_X1 output57 (.A(net57),
    .Z(result_o[17]));
 BUF_X1 output58 (.A(net58),
    .Z(result_o[18]));
 BUF_X1 output59 (.A(net59),
    .Z(result_o[19]));
 BUF_X1 output60 (.A(net60),
    .Z(result_o[1]));
 BUF_X1 output61 (.A(net61),
    .Z(result_o[20]));
 BUF_X1 output62 (.A(net62),
    .Z(result_o[21]));
 BUF_X1 output63 (.A(net63),
    .Z(result_o[22]));
 BUF_X1 output64 (.A(net64),
    .Z(result_o[23]));
 BUF_X1 output65 (.A(net65),
    .Z(result_o[24]));
 BUF_X1 output66 (.A(net66),
    .Z(result_o[25]));
 BUF_X1 output67 (.A(net67),
    .Z(result_o[26]));
 BUF_X1 output68 (.A(net68),
    .Z(result_o[27]));
 BUF_X1 output69 (.A(net69),
    .Z(result_o[28]));
 BUF_X1 output70 (.A(net70),
    .Z(result_o[29]));
 BUF_X1 output71 (.A(net71),
    .Z(result_o[2]));
 BUF_X1 output72 (.A(net72),
    .Z(result_o[30]));
 BUF_X1 output73 (.A(net73),
    .Z(result_o[31]));
 BUF_X1 output74 (.A(net74),
    .Z(result_o[3]));
 BUF_X1 output75 (.A(net75),
    .Z(result_o[4]));
 BUF_X1 output76 (.A(net76),
    .Z(result_o[5]));
 BUF_X1 output77 (.A(net77),
    .Z(result_o[6]));
 BUF_X1 output78 (.A(net78),
    .Z(result_o[7]));
 BUF_X1 output79 (.A(net79),
    .Z(result_o[8]));
 BUF_X1 output80 (.A(net80),
    .Z(result_o[9]));
 BUF_X4 max_cap81 (.A(_0247_),
    .Z(net81));
 BUF_X4 max_cap82 (.A(net83),
    .Z(net82));
 BUF_X4 max_cap83 (.A(_2120_),
    .Z(net83));
 BUF_X4 max_cap84 (.A(_2120_),
    .Z(net84));
 BUF_X4 max_cap85 (.A(net86),
    .Z(net85));
 CLKBUF_X3 max_cap86 (.A(net115),
    .Z(net86));
 BUF_X4 max_cap87 (.A(net115),
    .Z(net87));
 CLKBUF_X3 max_cap88 (.A(_2363_),
    .Z(net88));
 BUF_X8 max_cap89 (.A(net97),
    .Z(net89));
 BUF_X16 max_cap90 (.A(net131),
    .Z(net90));
 BUF_X4 max_cap91 (.A(net92),
    .Z(net91));
 BUF_X4 max_cap92 (.A(net93),
    .Z(net92));
 BUF_X4 max_cap93 (.A(net94),
    .Z(net93));
 CLKBUF_X3 wire94 (.A(net95),
    .Z(net94));
 CLKBUF_X3 max_cap95 (.A(_2269_),
    .Z(net95));
 BUF_X4 max_cap96 (.A(net125),
    .Z(net96));
 BUF_X1 rebuffer1 (.A(_1575_),
    .Z(net97));
 CLKBUF_X1 rebuffer2 (.A(net97),
    .Z(net98));
 BUF_X2 rebuffer3 (.A(_2127_),
    .Z(net99));
 CLKBUF_X1 rebuffer4 (.A(net99),
    .Z(net100));
 BUF_X8 split5 (.A(net109),
    .Z(net101));
 CLKBUF_X1 rebuffer6 (.A(_1546_),
    .Z(net102));
 BUF_X2 rebuffer7 (.A(net102),
    .Z(net103));
 BUF_X4 split8 (.A(net117),
    .Z(net104));
 CLKBUF_X3 split9 (.A(_1553_),
    .Z(net105));
 CLKBUF_X1 rebuffer10 (.A(_2051_),
    .Z(net106));
 CLKBUF_X1 rebuffer11 (.A(net106),
    .Z(net107));
 CLKBUF_X1 rebuffer12 (.A(_2214_),
    .Z(net108));
 BUF_X4 split13 (.A(_1549_),
    .Z(net109));
 CLKBUF_X2 split14 (.A(_1546_),
    .Z(net110));
 BUF_X2 split15 (.A(_1553_),
    .Z(net111));
 BUF_X4 rebuffer16 (.A(_1542_),
    .Z(net112));
 CLKBUF_X1 rebuffer17 (.A(_1542_),
    .Z(net113));
 BUF_X2 rebuffer18 (.A(_0232_),
    .Z(net114));
 BUF_X4 rebuffer19 (.A(_2114_),
    .Z(net115));
 BUF_X2 split20 (.A(_1505_),
    .Z(net116));
 BUF_X2 split21 (.A(_0232_),
    .Z(net117));
 BUF_X2 split22 (.A(_1542_),
    .Z(net118));
 CLKBUF_X1 rebuffer23 (.A(_2028_),
    .Z(net119));
 BUF_X8 split24 (.A(_0267_),
    .Z(net120));
 BUF_X1 split25 (.A(_1505_),
    .Z(net121));
 CLKBUF_X1 rebuffer26 (.A(net135),
    .Z(net122));
 CLKBUF_X1 rebuffer27 (.A(_1549_),
    .Z(net123));
 CLKBUF_X1 rebuffer28 (.A(_1549_),
    .Z(net124));
 CLKBUF_X1 rebuffer29 (.A(_2229_),
    .Z(net125));
 CLKBUF_X1 rebuffer30 (.A(net125),
    .Z(net126));
 BUF_X4 split31 (.A(net147),
    .Z(net127));
 CLKBUF_X3 split32 (.A(net134),
    .Z(net128));
 CLKBUF_X3 split33 (.A(_1620_),
    .Z(net129));
 CLKBUF_X1 rebuffer34 (.A(_2016_),
    .Z(net130));
 BUF_X2 rebuffer35 (.A(_1542_),
    .Z(net131));
 BUF_X8 split36 (.A(_0267_),
    .Z(net132));
 BUF_X2 rebuffer37 (.A(_1347_),
    .Z(net133));
 BUF_X4 split38 (.A(_1244_),
    .Z(net134));
 BUF_X4 rebuffer39 (.A(_1242_),
    .Z(net135));
 CLKBUF_X1 rebuffer40 (.A(_2373_),
    .Z(net136));
 CLKBUF_X1 rebuffer41 (.A(_1564_),
    .Z(net137));
 CLKBUF_X1 rebuffer42 (.A(_1564_),
    .Z(net138));
 CLKBUF_X1 rebuffer43 (.A(_2370_),
    .Z(net139));
 BUF_X2 rebuffer44 (.A(_1310_),
    .Z(net140));
 BUF_X1 rebuffer45 (.A(_2372_),
    .Z(net141));
 CLKBUF_X1 rebuffer46 (.A(net141),
    .Z(net142));
 BUF_X1 rebuffer47 (.A(net141),
    .Z(net143));
 BUF_X1 rebuffer48 (.A(net141),
    .Z(net144));
 CLKBUF_X1 rebuffer49 (.A(_1620_),
    .Z(net145));
 BUF_X4 rebuffer50 (.A(_1976_),
    .Z(net146));
 CLKBUF_X3 split51 (.A(net150),
    .Z(net147));
 CLKBUF_X1 rebuffer52 (.A(_1487_),
    .Z(net148));
 BUF_X2 rebuffer53 (.A(_2220_),
    .Z(net149));
 BUF_X1 split54 (.A(_0229_),
    .Z(net150));
 BUF_X4 split86 (.A(_1017_),
    .Z(net182));
 CLKBUF_X2 split91 (.A(_1017_),
    .Z(net187));
 BUF_X4 split96 (.A(_1018_),
    .Z(net192));
 CLKBUF_X3 split97 (.A(_1018_),
    .Z(net193));
 FILLCELL_X32 FILLER_0_0_1 ();
 FILLCELL_X32 FILLER_0_0_33 ();
 FILLCELL_X32 FILLER_0_0_65 ();
 FILLCELL_X32 FILLER_0_0_97 ();
 FILLCELL_X4 FILLER_0_0_129 ();
 FILLCELL_X4 FILLER_0_0_136 ();
 FILLCELL_X2 FILLER_0_0_140 ();
 FILLCELL_X1 FILLER_0_0_142 ();
 FILLCELL_X8 FILLER_0_0_146 ();
 FILLCELL_X1 FILLER_0_0_180 ();
 FILLCELL_X2 FILLER_0_0_197 ();
 FILLCELL_X1 FILLER_0_0_203 ();
 FILLCELL_X2 FILLER_0_0_220 ();
 FILLCELL_X1 FILLER_0_0_257 ();
 FILLCELL_X2 FILLER_0_0_285 ();
 FILLCELL_X32 FILLER_0_0_290 ();
 FILLCELL_X32 FILLER_0_0_322 ();
 FILLCELL_X32 FILLER_0_0_354 ();
 FILLCELL_X16 FILLER_0_0_386 ();
 FILLCELL_X4 FILLER_0_0_402 ();
 FILLCELL_X2 FILLER_0_0_406 ();
 FILLCELL_X32 FILLER_0_1_1 ();
 FILLCELL_X32 FILLER_0_1_33 ();
 FILLCELL_X32 FILLER_0_1_65 ();
 FILLCELL_X32 FILLER_0_1_97 ();
 FILLCELL_X16 FILLER_0_1_129 ();
 FILLCELL_X8 FILLER_0_1_145 ();
 FILLCELL_X4 FILLER_0_1_153 ();
 FILLCELL_X2 FILLER_0_1_157 ();
 FILLCELL_X1 FILLER_0_1_169 ();
 FILLCELL_X1 FILLER_0_1_205 ();
 FILLCELL_X1 FILLER_0_1_250 ();
 FILLCELL_X2 FILLER_0_1_287 ();
 FILLCELL_X32 FILLER_0_1_292 ();
 FILLCELL_X32 FILLER_0_1_324 ();
 FILLCELL_X32 FILLER_0_1_356 ();
 FILLCELL_X16 FILLER_0_1_388 ();
 FILLCELL_X4 FILLER_0_1_404 ();
 FILLCELL_X32 FILLER_0_2_1 ();
 FILLCELL_X32 FILLER_0_2_33 ();
 FILLCELL_X32 FILLER_0_2_65 ();
 FILLCELL_X32 FILLER_0_2_97 ();
 FILLCELL_X8 FILLER_0_2_129 ();
 FILLCELL_X4 FILLER_0_2_137 ();
 FILLCELL_X2 FILLER_0_2_141 ();
 FILLCELL_X2 FILLER_0_2_148 ();
 FILLCELL_X1 FILLER_0_2_150 ();
 FILLCELL_X2 FILLER_0_2_181 ();
 FILLCELL_X1 FILLER_0_2_199 ();
 FILLCELL_X2 FILLER_0_2_218 ();
 FILLCELL_X1 FILLER_0_2_232 ();
 FILLCELL_X8 FILLER_0_2_280 ();
 FILLCELL_X4 FILLER_0_2_288 ();
 FILLCELL_X1 FILLER_0_2_292 ();
 FILLCELL_X1 FILLER_0_2_305 ();
 FILLCELL_X32 FILLER_0_2_316 ();
 FILLCELL_X32 FILLER_0_2_348 ();
 FILLCELL_X16 FILLER_0_2_380 ();
 FILLCELL_X8 FILLER_0_2_396 ();
 FILLCELL_X4 FILLER_0_2_404 ();
 FILLCELL_X32 FILLER_0_3_1 ();
 FILLCELL_X8 FILLER_0_3_33 ();
 FILLCELL_X4 FILLER_0_3_41 ();
 FILLCELL_X4 FILLER_0_3_47 ();
 FILLCELL_X1 FILLER_0_3_51 ();
 FILLCELL_X8 FILLER_0_3_55 ();
 FILLCELL_X1 FILLER_0_3_63 ();
 FILLCELL_X32 FILLER_0_3_66 ();
 FILLCELL_X32 FILLER_0_3_98 ();
 FILLCELL_X4 FILLER_0_3_130 ();
 FILLCELL_X8 FILLER_0_3_148 ();
 FILLCELL_X4 FILLER_0_3_156 ();
 FILLCELL_X2 FILLER_0_3_160 ();
 FILLCELL_X1 FILLER_0_3_162 ();
 FILLCELL_X1 FILLER_0_3_186 ();
 FILLCELL_X2 FILLER_0_3_194 ();
 FILLCELL_X1 FILLER_0_3_211 ();
 FILLCELL_X1 FILLER_0_3_215 ();
 FILLCELL_X2 FILLER_0_3_220 ();
 FILLCELL_X1 FILLER_0_3_222 ();
 FILLCELL_X2 FILLER_0_3_234 ();
 FILLCELL_X1 FILLER_0_3_236 ();
 FILLCELL_X1 FILLER_0_3_243 ();
 FILLCELL_X8 FILLER_0_3_272 ();
 FILLCELL_X2 FILLER_0_3_280 ();
 FILLCELL_X1 FILLER_0_3_284 ();
 FILLCELL_X2 FILLER_0_3_297 ();
 FILLCELL_X8 FILLER_0_3_305 ();
 FILLCELL_X32 FILLER_0_3_315 ();
 FILLCELL_X32 FILLER_0_3_347 ();
 FILLCELL_X16 FILLER_0_3_379 ();
 FILLCELL_X8 FILLER_0_3_395 ();
 FILLCELL_X4 FILLER_0_3_403 ();
 FILLCELL_X1 FILLER_0_3_407 ();
 FILLCELL_X16 FILLER_0_4_1 ();
 FILLCELL_X1 FILLER_0_4_30 ();
 FILLCELL_X2 FILLER_0_4_34 ();
 FILLCELL_X32 FILLER_0_4_81 ();
 FILLCELL_X8 FILLER_0_4_113 ();
 FILLCELL_X4 FILLER_0_4_121 ();
 FILLCELL_X1 FILLER_0_4_125 ();
 FILLCELL_X1 FILLER_0_4_130 ();
 FILLCELL_X2 FILLER_0_4_144 ();
 FILLCELL_X1 FILLER_0_4_146 ();
 FILLCELL_X2 FILLER_0_4_150 ();
 FILLCELL_X1 FILLER_0_4_163 ();
 FILLCELL_X2 FILLER_0_4_177 ();
 FILLCELL_X2 FILLER_0_4_204 ();
 FILLCELL_X1 FILLER_0_4_213 ();
 FILLCELL_X4 FILLER_0_4_242 ();
 FILLCELL_X1 FILLER_0_4_246 ();
 FILLCELL_X1 FILLER_0_4_258 ();
 FILLCELL_X1 FILLER_0_4_261 ();
 FILLCELL_X1 FILLER_0_4_279 ();
 FILLCELL_X1 FILLER_0_4_288 ();
 FILLCELL_X8 FILLER_0_4_292 ();
 FILLCELL_X1 FILLER_0_4_310 ();
 FILLCELL_X32 FILLER_0_4_313 ();
 FILLCELL_X32 FILLER_0_4_345 ();
 FILLCELL_X16 FILLER_0_4_377 ();
 FILLCELL_X8 FILLER_0_4_393 ();
 FILLCELL_X4 FILLER_0_4_401 ();
 FILLCELL_X2 FILLER_0_4_405 ();
 FILLCELL_X1 FILLER_0_4_407 ();
 FILLCELL_X4 FILLER_0_5_1 ();
 FILLCELL_X2 FILLER_0_5_5 ();
 FILLCELL_X4 FILLER_0_5_10 ();
 FILLCELL_X2 FILLER_0_5_14 ();
 FILLCELL_X1 FILLER_0_5_39 ();
 FILLCELL_X1 FILLER_0_5_66 ();
 FILLCELL_X8 FILLER_0_5_101 ();
 FILLCELL_X1 FILLER_0_5_109 ();
 FILLCELL_X4 FILLER_0_5_113 ();
 FILLCELL_X2 FILLER_0_5_117 ();
 FILLCELL_X1 FILLER_0_5_119 ();
 FILLCELL_X2 FILLER_0_5_123 ();
 FILLCELL_X1 FILLER_0_5_125 ();
 FILLCELL_X1 FILLER_0_5_130 ();
 FILLCELL_X4 FILLER_0_5_147 ();
 FILLCELL_X1 FILLER_0_5_161 ();
 FILLCELL_X2 FILLER_0_5_165 ();
 FILLCELL_X2 FILLER_0_5_170 ();
 FILLCELL_X2 FILLER_0_5_176 ();
 FILLCELL_X1 FILLER_0_5_189 ();
 FILLCELL_X1 FILLER_0_5_195 ();
 FILLCELL_X1 FILLER_0_5_200 ();
 FILLCELL_X2 FILLER_0_5_203 ();
 FILLCELL_X2 FILLER_0_5_208 ();
 FILLCELL_X1 FILLER_0_5_210 ();
 FILLCELL_X4 FILLER_0_5_214 ();
 FILLCELL_X2 FILLER_0_5_232 ();
 FILLCELL_X1 FILLER_0_5_234 ();
 FILLCELL_X4 FILLER_0_5_241 ();
 FILLCELL_X2 FILLER_0_5_245 ();
 FILLCELL_X2 FILLER_0_5_257 ();
 FILLCELL_X2 FILLER_0_5_299 ();
 FILLCELL_X32 FILLER_0_5_317 ();
 FILLCELL_X32 FILLER_0_5_349 ();
 FILLCELL_X16 FILLER_0_5_381 ();
 FILLCELL_X8 FILLER_0_5_397 ();
 FILLCELL_X2 FILLER_0_5_405 ();
 FILLCELL_X1 FILLER_0_5_407 ();
 FILLCELL_X4 FILLER_0_6_1 ();
 FILLCELL_X1 FILLER_0_6_10 ();
 FILLCELL_X1 FILLER_0_6_29 ();
 FILLCELL_X2 FILLER_0_6_37 ();
 FILLCELL_X1 FILLER_0_6_46 ();
 FILLCELL_X2 FILLER_0_6_66 ();
 FILLCELL_X1 FILLER_0_6_68 ();
 FILLCELL_X2 FILLER_0_6_82 ();
 FILLCELL_X1 FILLER_0_6_84 ();
 FILLCELL_X1 FILLER_0_6_99 ();
 FILLCELL_X2 FILLER_0_6_108 ();
 FILLCELL_X1 FILLER_0_6_110 ();
 FILLCELL_X16 FILLER_0_6_153 ();
 FILLCELL_X4 FILLER_0_6_169 ();
 FILLCELL_X2 FILLER_0_6_173 ();
 FILLCELL_X2 FILLER_0_6_177 ();
 FILLCELL_X1 FILLER_0_6_179 ();
 FILLCELL_X4 FILLER_0_6_182 ();
 FILLCELL_X1 FILLER_0_6_192 ();
 FILLCELL_X1 FILLER_0_6_199 ();
 FILLCELL_X1 FILLER_0_6_204 ();
 FILLCELL_X1 FILLER_0_6_209 ();
 FILLCELL_X1 FILLER_0_6_214 ();
 FILLCELL_X1 FILLER_0_6_223 ();
 FILLCELL_X1 FILLER_0_6_265 ();
 FILLCELL_X4 FILLER_0_6_289 ();
 FILLCELL_X1 FILLER_0_6_293 ();
 FILLCELL_X1 FILLER_0_6_306 ();
 FILLCELL_X32 FILLER_0_6_322 ();
 FILLCELL_X32 FILLER_0_6_354 ();
 FILLCELL_X16 FILLER_0_6_386 ();
 FILLCELL_X4 FILLER_0_6_402 ();
 FILLCELL_X2 FILLER_0_6_406 ();
 FILLCELL_X4 FILLER_0_7_1 ();
 FILLCELL_X1 FILLER_0_7_5 ();
 FILLCELL_X1 FILLER_0_7_18 ();
 FILLCELL_X1 FILLER_0_7_27 ();
 FILLCELL_X1 FILLER_0_7_38 ();
 FILLCELL_X1 FILLER_0_7_50 ();
 FILLCELL_X2 FILLER_0_7_57 ();
 FILLCELL_X1 FILLER_0_7_59 ();
 FILLCELL_X2 FILLER_0_7_68 ();
 FILLCELL_X1 FILLER_0_7_70 ();
 FILLCELL_X1 FILLER_0_7_75 ();
 FILLCELL_X4 FILLER_0_7_81 ();
 FILLCELL_X4 FILLER_0_7_133 ();
 FILLCELL_X1 FILLER_0_7_137 ();
 FILLCELL_X1 FILLER_0_7_154 ();
 FILLCELL_X1 FILLER_0_7_162 ();
 FILLCELL_X2 FILLER_0_7_165 ();
 FILLCELL_X1 FILLER_0_7_180 ();
 FILLCELL_X8 FILLER_0_7_189 ();
 FILLCELL_X4 FILLER_0_7_197 ();
 FILLCELL_X2 FILLER_0_7_201 ();
 FILLCELL_X1 FILLER_0_7_203 ();
 FILLCELL_X4 FILLER_0_7_211 ();
 FILLCELL_X2 FILLER_0_7_215 ();
 FILLCELL_X1 FILLER_0_7_217 ();
 FILLCELL_X2 FILLER_0_7_223 ();
 FILLCELL_X1 FILLER_0_7_232 ();
 FILLCELL_X16 FILLER_0_7_236 ();
 FILLCELL_X2 FILLER_0_7_252 ();
 FILLCELL_X8 FILLER_0_7_261 ();
 FILLCELL_X2 FILLER_0_7_269 ();
 FILLCELL_X1 FILLER_0_7_271 ();
 FILLCELL_X1 FILLER_0_7_276 ();
 FILLCELL_X1 FILLER_0_7_299 ();
 FILLCELL_X1 FILLER_0_7_313 ();
 FILLCELL_X32 FILLER_0_7_317 ();
 FILLCELL_X32 FILLER_0_7_349 ();
 FILLCELL_X16 FILLER_0_7_381 ();
 FILLCELL_X8 FILLER_0_7_397 ();
 FILLCELL_X2 FILLER_0_7_405 ();
 FILLCELL_X1 FILLER_0_7_407 ();
 FILLCELL_X2 FILLER_0_8_14 ();
 FILLCELL_X2 FILLER_0_8_43 ();
 FILLCELL_X8 FILLER_0_8_48 ();
 FILLCELL_X4 FILLER_0_8_56 ();
 FILLCELL_X2 FILLER_0_8_60 ();
 FILLCELL_X1 FILLER_0_8_77 ();
 FILLCELL_X8 FILLER_0_8_81 ();
 FILLCELL_X4 FILLER_0_8_89 ();
 FILLCELL_X4 FILLER_0_8_97 ();
 FILLCELL_X8 FILLER_0_8_138 ();
 FILLCELL_X1 FILLER_0_8_146 ();
 FILLCELL_X2 FILLER_0_8_149 ();
 FILLCELL_X16 FILLER_0_8_154 ();
 FILLCELL_X4 FILLER_0_8_170 ();
 FILLCELL_X1 FILLER_0_8_177 ();
 FILLCELL_X2 FILLER_0_8_189 ();
 FILLCELL_X4 FILLER_0_8_200 ();
 FILLCELL_X16 FILLER_0_8_210 ();
 FILLCELL_X2 FILLER_0_8_226 ();
 FILLCELL_X1 FILLER_0_8_228 ();
 FILLCELL_X1 FILLER_0_8_236 ();
 FILLCELL_X8 FILLER_0_8_239 ();
 FILLCELL_X4 FILLER_0_8_257 ();
 FILLCELL_X2 FILLER_0_8_261 ();
 FILLCELL_X2 FILLER_0_8_268 ();
 FILLCELL_X4 FILLER_0_8_273 ();
 FILLCELL_X1 FILLER_0_8_277 ();
 FILLCELL_X1 FILLER_0_8_280 ();
 FILLCELL_X1 FILLER_0_8_291 ();
 FILLCELL_X1 FILLER_0_8_294 ();
 FILLCELL_X1 FILLER_0_8_301 ();
 FILLCELL_X2 FILLER_0_8_310 ();
 FILLCELL_X1 FILLER_0_8_312 ();
 FILLCELL_X32 FILLER_0_8_325 ();
 FILLCELL_X32 FILLER_0_8_357 ();
 FILLCELL_X16 FILLER_0_8_389 ();
 FILLCELL_X2 FILLER_0_8_405 ();
 FILLCELL_X1 FILLER_0_8_407 ();
 FILLCELL_X4 FILLER_0_9_1 ();
 FILLCELL_X2 FILLER_0_9_5 ();
 FILLCELL_X4 FILLER_0_9_21 ();
 FILLCELL_X2 FILLER_0_9_25 ();
 FILLCELL_X2 FILLER_0_9_34 ();
 FILLCELL_X1 FILLER_0_9_36 ();
 FILLCELL_X2 FILLER_0_9_44 ();
 FILLCELL_X1 FILLER_0_9_49 ();
 FILLCELL_X1 FILLER_0_9_54 ();
 FILLCELL_X2 FILLER_0_9_69 ();
 FILLCELL_X1 FILLER_0_9_83 ();
 FILLCELL_X2 FILLER_0_9_89 ();
 FILLCELL_X1 FILLER_0_9_91 ();
 FILLCELL_X2 FILLER_0_9_99 ();
 FILLCELL_X1 FILLER_0_9_141 ();
 FILLCELL_X1 FILLER_0_9_146 ();
 FILLCELL_X4 FILLER_0_9_151 ();
 FILLCELL_X8 FILLER_0_9_159 ();
 FILLCELL_X1 FILLER_0_9_167 ();
 FILLCELL_X2 FILLER_0_9_171 ();
 FILLCELL_X2 FILLER_0_9_213 ();
 FILLCELL_X1 FILLER_0_9_215 ();
 FILLCELL_X1 FILLER_0_9_227 ();
 FILLCELL_X32 FILLER_0_9_323 ();
 FILLCELL_X32 FILLER_0_9_355 ();
 FILLCELL_X16 FILLER_0_9_387 ();
 FILLCELL_X4 FILLER_0_9_403 ();
 FILLCELL_X1 FILLER_0_9_407 ();
 FILLCELL_X4 FILLER_0_10_1 ();
 FILLCELL_X1 FILLER_0_10_5 ();
 FILLCELL_X8 FILLER_0_10_22 ();
 FILLCELL_X2 FILLER_0_10_30 ();
 FILLCELL_X1 FILLER_0_10_40 ();
 FILLCELL_X1 FILLER_0_10_58 ();
 FILLCELL_X4 FILLER_0_10_73 ();
 FILLCELL_X1 FILLER_0_10_77 ();
 FILLCELL_X4 FILLER_0_10_81 ();
 FILLCELL_X1 FILLER_0_10_88 ();
 FILLCELL_X1 FILLER_0_10_92 ();
 FILLCELL_X1 FILLER_0_10_95 ();
 FILLCELL_X1 FILLER_0_10_135 ();
 FILLCELL_X1 FILLER_0_10_139 ();
 FILLCELL_X2 FILLER_0_10_153 ();
 FILLCELL_X1 FILLER_0_10_165 ();
 FILLCELL_X2 FILLER_0_10_173 ();
 FILLCELL_X2 FILLER_0_10_178 ();
 FILLCELL_X2 FILLER_0_10_192 ();
 FILLCELL_X1 FILLER_0_10_196 ();
 FILLCELL_X8 FILLER_0_10_200 ();
 FILLCELL_X1 FILLER_0_10_208 ();
 FILLCELL_X1 FILLER_0_10_213 ();
 FILLCELL_X4 FILLER_0_10_217 ();
 FILLCELL_X1 FILLER_0_10_221 ();
 FILLCELL_X16 FILLER_0_10_242 ();
 FILLCELL_X4 FILLER_0_10_258 ();
 FILLCELL_X2 FILLER_0_10_262 ();
 FILLCELL_X1 FILLER_0_10_264 ();
 FILLCELL_X4 FILLER_0_10_268 ();
 FILLCELL_X1 FILLER_0_10_272 ();
 FILLCELL_X4 FILLER_0_10_275 ();
 FILLCELL_X2 FILLER_0_10_279 ();
 FILLCELL_X1 FILLER_0_10_281 ();
 FILLCELL_X4 FILLER_0_10_293 ();
 FILLCELL_X32 FILLER_0_10_324 ();
 FILLCELL_X32 FILLER_0_10_356 ();
 FILLCELL_X16 FILLER_0_10_388 ();
 FILLCELL_X4 FILLER_0_10_404 ();
 FILLCELL_X4 FILLER_0_11_1 ();
 FILLCELL_X2 FILLER_0_11_5 ();
 FILLCELL_X1 FILLER_0_11_25 ();
 FILLCELL_X2 FILLER_0_11_38 ();
 FILLCELL_X4 FILLER_0_11_47 ();
 FILLCELL_X2 FILLER_0_11_51 ();
 FILLCELL_X1 FILLER_0_11_53 ();
 FILLCELL_X2 FILLER_0_11_63 ();
 FILLCELL_X8 FILLER_0_11_68 ();
 FILLCELL_X1 FILLER_0_11_76 ();
 FILLCELL_X1 FILLER_0_11_79 ();
 FILLCELL_X4 FILLER_0_11_84 ();
 FILLCELL_X1 FILLER_0_11_88 ();
 FILLCELL_X4 FILLER_0_11_93 ();
 FILLCELL_X2 FILLER_0_11_97 ();
 FILLCELL_X1 FILLER_0_11_99 ();
 FILLCELL_X1 FILLER_0_11_108 ();
 FILLCELL_X1 FILLER_0_11_112 ();
 FILLCELL_X1 FILLER_0_11_119 ();
 FILLCELL_X2 FILLER_0_11_131 ();
 FILLCELL_X8 FILLER_0_11_135 ();
 FILLCELL_X1 FILLER_0_11_143 ();
 FILLCELL_X4 FILLER_0_11_149 ();
 FILLCELL_X1 FILLER_0_11_153 ();
 FILLCELL_X4 FILLER_0_11_156 ();
 FILLCELL_X2 FILLER_0_11_165 ();
 FILLCELL_X1 FILLER_0_11_167 ();
 FILLCELL_X4 FILLER_0_11_172 ();
 FILLCELL_X4 FILLER_0_11_180 ();
 FILLCELL_X2 FILLER_0_11_184 ();
 FILLCELL_X1 FILLER_0_11_186 ();
 FILLCELL_X8 FILLER_0_11_191 ();
 FILLCELL_X2 FILLER_0_11_206 ();
 FILLCELL_X4 FILLER_0_11_210 ();
 FILLCELL_X1 FILLER_0_11_214 ();
 FILLCELL_X2 FILLER_0_11_220 ();
 FILLCELL_X1 FILLER_0_11_222 ();
 FILLCELL_X4 FILLER_0_11_227 ();
 FILLCELL_X2 FILLER_0_11_231 ();
 FILLCELL_X1 FILLER_0_11_233 ();
 FILLCELL_X1 FILLER_0_11_240 ();
 FILLCELL_X16 FILLER_0_11_243 ();
 FILLCELL_X8 FILLER_0_11_259 ();
 FILLCELL_X4 FILLER_0_11_267 ();
 FILLCELL_X2 FILLER_0_11_271 ();
 FILLCELL_X1 FILLER_0_11_285 ();
 FILLCELL_X1 FILLER_0_11_308 ();
 FILLCELL_X32 FILLER_0_11_332 ();
 FILLCELL_X32 FILLER_0_11_364 ();
 FILLCELL_X8 FILLER_0_11_396 ();
 FILLCELL_X4 FILLER_0_11_404 ();
 FILLCELL_X16 FILLER_0_12_1 ();
 FILLCELL_X4 FILLER_0_12_31 ();
 FILLCELL_X2 FILLER_0_12_35 ();
 FILLCELL_X1 FILLER_0_12_37 ();
 FILLCELL_X16 FILLER_0_12_40 ();
 FILLCELL_X2 FILLER_0_12_89 ();
 FILLCELL_X1 FILLER_0_12_91 ();
 FILLCELL_X8 FILLER_0_12_99 ();
 FILLCELL_X1 FILLER_0_12_107 ();
 FILLCELL_X1 FILLER_0_12_110 ();
 FILLCELL_X1 FILLER_0_12_118 ();
 FILLCELL_X2 FILLER_0_12_132 ();
 FILLCELL_X2 FILLER_0_12_146 ();
 FILLCELL_X8 FILLER_0_12_157 ();
 FILLCELL_X4 FILLER_0_12_165 ();
 FILLCELL_X2 FILLER_0_12_169 ();
 FILLCELL_X2 FILLER_0_12_197 ();
 FILLCELL_X1 FILLER_0_12_199 ();
 FILLCELL_X1 FILLER_0_12_218 ();
 FILLCELL_X1 FILLER_0_12_221 ();
 FILLCELL_X2 FILLER_0_12_232 ();
 FILLCELL_X1 FILLER_0_12_234 ();
 FILLCELL_X4 FILLER_0_12_241 ();
 FILLCELL_X1 FILLER_0_12_245 ();
 FILLCELL_X2 FILLER_0_12_257 ();
 FILLCELL_X1 FILLER_0_12_277 ();
 FILLCELL_X2 FILLER_0_12_296 ();
 FILLCELL_X1 FILLER_0_12_301 ();
 FILLCELL_X32 FILLER_0_12_335 ();
 FILLCELL_X32 FILLER_0_12_367 ();
 FILLCELL_X8 FILLER_0_12_399 ();
 FILLCELL_X1 FILLER_0_12_407 ();
 FILLCELL_X16 FILLER_0_13_1 ();
 FILLCELL_X2 FILLER_0_13_17 ();
 FILLCELL_X1 FILLER_0_13_19 ();
 FILLCELL_X4 FILLER_0_13_29 ();
 FILLCELL_X1 FILLER_0_13_51 ();
 FILLCELL_X8 FILLER_0_13_68 ();
 FILLCELL_X4 FILLER_0_13_76 ();
 FILLCELL_X1 FILLER_0_13_80 ();
 FILLCELL_X4 FILLER_0_13_83 ();
 FILLCELL_X8 FILLER_0_13_89 ();
 FILLCELL_X2 FILLER_0_13_97 ();
 FILLCELL_X1 FILLER_0_13_99 ();
 FILLCELL_X4 FILLER_0_13_103 ();
 FILLCELL_X1 FILLER_0_13_107 ();
 FILLCELL_X2 FILLER_0_13_114 ();
 FILLCELL_X1 FILLER_0_13_116 ();
 FILLCELL_X2 FILLER_0_13_119 ();
 FILLCELL_X4 FILLER_0_13_133 ();
 FILLCELL_X2 FILLER_0_13_137 ();
 FILLCELL_X1 FILLER_0_13_154 ();
 FILLCELL_X4 FILLER_0_13_181 ();
 FILLCELL_X2 FILLER_0_13_185 ();
 FILLCELL_X1 FILLER_0_13_187 ();
 FILLCELL_X2 FILLER_0_13_200 ();
 FILLCELL_X1 FILLER_0_13_202 ();
 FILLCELL_X8 FILLER_0_13_236 ();
 FILLCELL_X4 FILLER_0_13_244 ();
 FILLCELL_X1 FILLER_0_13_248 ();
 FILLCELL_X4 FILLER_0_13_259 ();
 FILLCELL_X2 FILLER_0_13_263 ();
 FILLCELL_X1 FILLER_0_13_265 ();
 FILLCELL_X1 FILLER_0_13_275 ();
 FILLCELL_X2 FILLER_0_13_282 ();
 FILLCELL_X32 FILLER_0_13_318 ();
 FILLCELL_X32 FILLER_0_13_350 ();
 FILLCELL_X16 FILLER_0_13_382 ();
 FILLCELL_X8 FILLER_0_13_398 ();
 FILLCELL_X2 FILLER_0_13_406 ();
 FILLCELL_X8 FILLER_0_14_1 ();
 FILLCELL_X1 FILLER_0_14_9 ();
 FILLCELL_X1 FILLER_0_14_17 ();
 FILLCELL_X8 FILLER_0_14_23 ();
 FILLCELL_X1 FILLER_0_14_31 ();
 FILLCELL_X2 FILLER_0_14_47 ();
 FILLCELL_X1 FILLER_0_14_64 ();
 FILLCELL_X1 FILLER_0_14_72 ();
 FILLCELL_X16 FILLER_0_14_80 ();
 FILLCELL_X2 FILLER_0_14_96 ();
 FILLCELL_X1 FILLER_0_14_111 ();
 FILLCELL_X2 FILLER_0_14_128 ();
 FILLCELL_X1 FILLER_0_14_130 ();
 FILLCELL_X8 FILLER_0_14_135 ();
 FILLCELL_X1 FILLER_0_14_143 ();
 FILLCELL_X2 FILLER_0_14_156 ();
 FILLCELL_X2 FILLER_0_14_161 ();
 FILLCELL_X2 FILLER_0_14_166 ();
 FILLCELL_X1 FILLER_0_14_180 ();
 FILLCELL_X4 FILLER_0_14_187 ();
 FILLCELL_X1 FILLER_0_14_191 ();
 FILLCELL_X4 FILLER_0_14_198 ();
 FILLCELL_X2 FILLER_0_14_202 ();
 FILLCELL_X1 FILLER_0_14_204 ();
 FILLCELL_X2 FILLER_0_14_214 ();
 FILLCELL_X1 FILLER_0_14_216 ();
 FILLCELL_X2 FILLER_0_14_224 ();
 FILLCELL_X1 FILLER_0_14_226 ();
 FILLCELL_X2 FILLER_0_14_231 ();
 FILLCELL_X2 FILLER_0_14_239 ();
 FILLCELL_X4 FILLER_0_14_246 ();
 FILLCELL_X2 FILLER_0_14_250 ();
 FILLCELL_X1 FILLER_0_14_268 ();
 FILLCELL_X4 FILLER_0_14_296 ();
 FILLCELL_X16 FILLER_0_14_309 ();
 FILLCELL_X8 FILLER_0_14_325 ();
 FILLCELL_X4 FILLER_0_14_333 ();
 FILLCELL_X1 FILLER_0_14_337 ();
 FILLCELL_X32 FILLER_0_14_340 ();
 FILLCELL_X32 FILLER_0_14_372 ();
 FILLCELL_X4 FILLER_0_14_404 ();
 FILLCELL_X8 FILLER_0_15_1 ();
 FILLCELL_X1 FILLER_0_15_26 ();
 FILLCELL_X1 FILLER_0_15_81 ();
 FILLCELL_X2 FILLER_0_15_107 ();
 FILLCELL_X1 FILLER_0_15_126 ();
 FILLCELL_X2 FILLER_0_15_131 ();
 FILLCELL_X1 FILLER_0_15_133 ();
 FILLCELL_X2 FILLER_0_15_136 ();
 FILLCELL_X1 FILLER_0_15_138 ();
 FILLCELL_X1 FILLER_0_15_142 ();
 FILLCELL_X2 FILLER_0_15_146 ();
 FILLCELL_X1 FILLER_0_15_148 ();
 FILLCELL_X4 FILLER_0_15_159 ();
 FILLCELL_X8 FILLER_0_15_172 ();
 FILLCELL_X2 FILLER_0_15_180 ();
 FILLCELL_X1 FILLER_0_15_192 ();
 FILLCELL_X4 FILLER_0_15_198 ();
 FILLCELL_X1 FILLER_0_15_202 ();
 FILLCELL_X2 FILLER_0_15_216 ();
 FILLCELL_X1 FILLER_0_15_218 ();
 FILLCELL_X2 FILLER_0_15_221 ();
 FILLCELL_X2 FILLER_0_15_229 ();
 FILLCELL_X8 FILLER_0_15_257 ();
 FILLCELL_X2 FILLER_0_15_265 ();
 FILLCELL_X1 FILLER_0_15_267 ();
 FILLCELL_X4 FILLER_0_15_298 ();
 FILLCELL_X1 FILLER_0_15_302 ();
 FILLCELL_X16 FILLER_0_15_306 ();
 FILLCELL_X8 FILLER_0_15_322 ();
 FILLCELL_X4 FILLER_0_15_330 ();
 FILLCELL_X2 FILLER_0_15_334 ();
 FILLCELL_X32 FILLER_0_15_346 ();
 FILLCELL_X16 FILLER_0_15_378 ();
 FILLCELL_X8 FILLER_0_15_394 ();
 FILLCELL_X4 FILLER_0_15_402 ();
 FILLCELL_X2 FILLER_0_15_406 ();
 FILLCELL_X8 FILLER_0_16_1 ();
 FILLCELL_X1 FILLER_0_16_9 ();
 FILLCELL_X16 FILLER_0_16_17 ();
 FILLCELL_X2 FILLER_0_16_33 ();
 FILLCELL_X1 FILLER_0_16_35 ();
 FILLCELL_X2 FILLER_0_16_48 ();
 FILLCELL_X1 FILLER_0_16_58 ();
 FILLCELL_X4 FILLER_0_16_67 ();
 FILLCELL_X4 FILLER_0_16_78 ();
 FILLCELL_X2 FILLER_0_16_86 ();
 FILLCELL_X4 FILLER_0_16_90 ();
 FILLCELL_X1 FILLER_0_16_94 ();
 FILLCELL_X1 FILLER_0_16_99 ();
 FILLCELL_X1 FILLER_0_16_118 ();
 FILLCELL_X8 FILLER_0_16_125 ();
 FILLCELL_X1 FILLER_0_16_139 ();
 FILLCELL_X4 FILLER_0_16_152 ();
 FILLCELL_X2 FILLER_0_16_156 ();
 FILLCELL_X2 FILLER_0_16_170 ();
 FILLCELL_X1 FILLER_0_16_172 ();
 FILLCELL_X2 FILLER_0_16_179 ();
 FILLCELL_X4 FILLER_0_16_190 ();
 FILLCELL_X1 FILLER_0_16_194 ();
 FILLCELL_X1 FILLER_0_16_207 ();
 FILLCELL_X4 FILLER_0_16_212 ();
 FILLCELL_X2 FILLER_0_16_216 ();
 FILLCELL_X1 FILLER_0_16_218 ();
 FILLCELL_X4 FILLER_0_16_235 ();
 FILLCELL_X8 FILLER_0_16_259 ();
 FILLCELL_X1 FILLER_0_16_303 ();
 FILLCELL_X4 FILLER_0_16_314 ();
 FILLCELL_X2 FILLER_0_16_318 ();
 FILLCELL_X2 FILLER_0_16_330 ();
 FILLCELL_X1 FILLER_0_16_332 ();
 FILLCELL_X2 FILLER_0_16_347 ();
 FILLCELL_X16 FILLER_0_16_355 ();
 FILLCELL_X8 FILLER_0_16_373 ();
 FILLCELL_X4 FILLER_0_16_381 ();
 FILLCELL_X2 FILLER_0_16_385 ();
 FILLCELL_X4 FILLER_0_16_389 ();
 FILLCELL_X2 FILLER_0_16_393 ();
 FILLCELL_X8 FILLER_0_16_397 ();
 FILLCELL_X2 FILLER_0_16_405 ();
 FILLCELL_X1 FILLER_0_16_407 ();
 FILLCELL_X8 FILLER_0_17_1 ();
 FILLCELL_X2 FILLER_0_17_9 ();
 FILLCELL_X8 FILLER_0_17_26 ();
 FILLCELL_X4 FILLER_0_17_34 ();
 FILLCELL_X2 FILLER_0_17_38 ();
 FILLCELL_X1 FILLER_0_17_40 ();
 FILLCELL_X2 FILLER_0_17_50 ();
 FILLCELL_X1 FILLER_0_17_55 ();
 FILLCELL_X8 FILLER_0_17_61 ();
 FILLCELL_X4 FILLER_0_17_69 ();
 FILLCELL_X1 FILLER_0_17_90 ();
 FILLCELL_X4 FILLER_0_17_102 ();
 FILLCELL_X1 FILLER_0_17_109 ();
 FILLCELL_X4 FILLER_0_17_116 ();
 FILLCELL_X2 FILLER_0_17_124 ();
 FILLCELL_X1 FILLER_0_17_126 ();
 FILLCELL_X1 FILLER_0_17_129 ();
 FILLCELL_X2 FILLER_0_17_140 ();
 FILLCELL_X1 FILLER_0_17_142 ();
 FILLCELL_X1 FILLER_0_17_151 ();
 FILLCELL_X1 FILLER_0_17_155 ();
 FILLCELL_X4 FILLER_0_17_159 ();
 FILLCELL_X1 FILLER_0_17_163 ();
 FILLCELL_X4 FILLER_0_17_169 ();
 FILLCELL_X8 FILLER_0_17_176 ();
 FILLCELL_X1 FILLER_0_17_184 ();
 FILLCELL_X16 FILLER_0_17_219 ();
 FILLCELL_X2 FILLER_0_17_235 ();
 FILLCELL_X8 FILLER_0_17_253 ();
 FILLCELL_X4 FILLER_0_17_261 ();
 FILLCELL_X1 FILLER_0_17_265 ();
 FILLCELL_X1 FILLER_0_17_278 ();
 FILLCELL_X1 FILLER_0_17_292 ();
 FILLCELL_X2 FILLER_0_17_297 ();
 FILLCELL_X1 FILLER_0_17_299 ();
 FILLCELL_X4 FILLER_0_17_302 ();
 FILLCELL_X1 FILLER_0_17_306 ();
 FILLCELL_X2 FILLER_0_17_336 ();
 FILLCELL_X1 FILLER_0_17_338 ();
 FILLCELL_X8 FILLER_0_17_341 ();
 FILLCELL_X2 FILLER_0_17_349 ();
 FILLCELL_X1 FILLER_0_17_378 ();
 FILLCELL_X8 FILLER_0_18_1 ();
 FILLCELL_X1 FILLER_0_18_9 ();
 FILLCELL_X1 FILLER_0_18_22 ();
 FILLCELL_X1 FILLER_0_18_26 ();
 FILLCELL_X1 FILLER_0_18_38 ();
 FILLCELL_X2 FILLER_0_18_45 ();
 FILLCELL_X1 FILLER_0_18_47 ();
 FILLCELL_X1 FILLER_0_18_65 ();
 FILLCELL_X1 FILLER_0_18_73 ();
 FILLCELL_X1 FILLER_0_18_78 ();
 FILLCELL_X1 FILLER_0_18_92 ();
 FILLCELL_X1 FILLER_0_18_111 ();
 FILLCELL_X16 FILLER_0_18_114 ();
 FILLCELL_X1 FILLER_0_18_134 ();
 FILLCELL_X1 FILLER_0_18_138 ();
 FILLCELL_X1 FILLER_0_18_141 ();
 FILLCELL_X1 FILLER_0_18_145 ();
 FILLCELL_X1 FILLER_0_18_184 ();
 FILLCELL_X8 FILLER_0_18_191 ();
 FILLCELL_X1 FILLER_0_18_199 ();
 FILLCELL_X16 FILLER_0_18_226 ();
 FILLCELL_X1 FILLER_0_18_242 ();
 FILLCELL_X1 FILLER_0_18_253 ();
 FILLCELL_X1 FILLER_0_18_259 ();
 FILLCELL_X4 FILLER_0_18_269 ();
 FILLCELL_X1 FILLER_0_18_273 ();
 FILLCELL_X2 FILLER_0_18_278 ();
 FILLCELL_X16 FILLER_0_18_282 ();
 FILLCELL_X8 FILLER_0_18_298 ();
 FILLCELL_X4 FILLER_0_18_306 ();
 FILLCELL_X2 FILLER_0_18_310 ();
 FILLCELL_X4 FILLER_0_18_337 ();
 FILLCELL_X4 FILLER_0_18_368 ();
 FILLCELL_X8 FILLER_0_19_1 ();
 FILLCELL_X4 FILLER_0_19_9 ();
 FILLCELL_X4 FILLER_0_19_26 ();
 FILLCELL_X2 FILLER_0_19_34 ();
 FILLCELL_X4 FILLER_0_19_51 ();
 FILLCELL_X2 FILLER_0_19_55 ();
 FILLCELL_X1 FILLER_0_19_57 ();
 FILLCELL_X1 FILLER_0_19_62 ();
 FILLCELL_X8 FILLER_0_19_70 ();
 FILLCELL_X4 FILLER_0_19_78 ();
 FILLCELL_X1 FILLER_0_19_82 ();
 FILLCELL_X1 FILLER_0_19_98 ();
 FILLCELL_X2 FILLER_0_19_106 ();
 FILLCELL_X1 FILLER_0_19_115 ();
 FILLCELL_X2 FILLER_0_19_122 ();
 FILLCELL_X1 FILLER_0_19_127 ();
 FILLCELL_X1 FILLER_0_19_135 ();
 FILLCELL_X1 FILLER_0_19_140 ();
 FILLCELL_X2 FILLER_0_19_149 ();
 FILLCELL_X8 FILLER_0_19_161 ();
 FILLCELL_X2 FILLER_0_19_169 ();
 FILLCELL_X2 FILLER_0_19_175 ();
 FILLCELL_X1 FILLER_0_19_177 ();
 FILLCELL_X1 FILLER_0_19_227 ();
 FILLCELL_X16 FILLER_0_19_230 ();
 FILLCELL_X1 FILLER_0_19_246 ();
 FILLCELL_X4 FILLER_0_19_279 ();
 FILLCELL_X8 FILLER_0_19_285 ();
 FILLCELL_X4 FILLER_0_19_293 ();
 FILLCELL_X2 FILLER_0_19_306 ();
 FILLCELL_X1 FILLER_0_19_308 ();
 FILLCELL_X1 FILLER_0_19_318 ();
 FILLCELL_X1 FILLER_0_19_322 ();
 FILLCELL_X1 FILLER_0_19_325 ();
 FILLCELL_X2 FILLER_0_19_336 ();
 FILLCELL_X2 FILLER_0_19_342 ();
 FILLCELL_X8 FILLER_0_19_346 ();
 FILLCELL_X2 FILLER_0_19_354 ();
 FILLCELL_X1 FILLER_0_19_356 ();
 FILLCELL_X4 FILLER_0_19_367 ();
 FILLCELL_X8 FILLER_0_19_374 ();
 FILLCELL_X1 FILLER_0_19_382 ();
 FILLCELL_X2 FILLER_0_19_403 ();
 FILLCELL_X16 FILLER_0_20_1 ();
 FILLCELL_X2 FILLER_0_20_17 ();
 FILLCELL_X16 FILLER_0_20_22 ();
 FILLCELL_X8 FILLER_0_20_38 ();
 FILLCELL_X1 FILLER_0_20_46 ();
 FILLCELL_X2 FILLER_0_20_62 ();
 FILLCELL_X2 FILLER_0_20_78 ();
 FILLCELL_X1 FILLER_0_20_80 ();
 FILLCELL_X1 FILLER_0_20_85 ();
 FILLCELL_X2 FILLER_0_20_93 ();
 FILLCELL_X1 FILLER_0_20_95 ();
 FILLCELL_X2 FILLER_0_20_100 ();
 FILLCELL_X1 FILLER_0_20_102 ();
 FILLCELL_X4 FILLER_0_20_108 ();
 FILLCELL_X2 FILLER_0_20_112 ();
 FILLCELL_X2 FILLER_0_20_127 ();
 FILLCELL_X4 FILLER_0_20_132 ();
 FILLCELL_X2 FILLER_0_20_136 ();
 FILLCELL_X4 FILLER_0_20_148 ();
 FILLCELL_X2 FILLER_0_20_152 ();
 FILLCELL_X1 FILLER_0_20_154 ();
 FILLCELL_X2 FILLER_0_20_167 ();
 FILLCELL_X2 FILLER_0_20_175 ();
 FILLCELL_X1 FILLER_0_20_179 ();
 FILLCELL_X2 FILLER_0_20_190 ();
 FILLCELL_X2 FILLER_0_20_221 ();
 FILLCELL_X1 FILLER_0_20_223 ();
 FILLCELL_X1 FILLER_0_20_230 ();
 FILLCELL_X1 FILLER_0_20_237 ();
 FILLCELL_X4 FILLER_0_20_240 ();
 FILLCELL_X2 FILLER_0_20_244 ();
 FILLCELL_X1 FILLER_0_20_246 ();
 FILLCELL_X4 FILLER_0_20_250 ();
 FILLCELL_X1 FILLER_0_20_254 ();
 FILLCELL_X2 FILLER_0_20_313 ();
 FILLCELL_X1 FILLER_0_20_315 ();
 FILLCELL_X4 FILLER_0_20_328 ();
 FILLCELL_X1 FILLER_0_20_332 ();
 FILLCELL_X16 FILLER_0_20_359 ();
 FILLCELL_X8 FILLER_0_20_375 ();
 FILLCELL_X1 FILLER_0_20_383 ();
 FILLCELL_X1 FILLER_0_20_404 ();
 FILLCELL_X16 FILLER_0_21_1 ();
 FILLCELL_X1 FILLER_0_21_17 ();
 FILLCELL_X8 FILLER_0_21_24 ();
 FILLCELL_X4 FILLER_0_21_32 ();
 FILLCELL_X2 FILLER_0_21_36 ();
 FILLCELL_X1 FILLER_0_21_38 ();
 FILLCELL_X8 FILLER_0_21_45 ();
 FILLCELL_X4 FILLER_0_21_53 ();
 FILLCELL_X2 FILLER_0_21_57 ();
 FILLCELL_X2 FILLER_0_21_67 ();
 FILLCELL_X1 FILLER_0_21_73 ();
 FILLCELL_X4 FILLER_0_21_77 ();
 FILLCELL_X2 FILLER_0_21_81 ();
 FILLCELL_X2 FILLER_0_21_94 ();
 FILLCELL_X4 FILLER_0_21_100 ();
 FILLCELL_X2 FILLER_0_21_104 ();
 FILLCELL_X4 FILLER_0_21_115 ();
 FILLCELL_X2 FILLER_0_21_119 ();
 FILLCELL_X4 FILLER_0_21_143 ();
 FILLCELL_X2 FILLER_0_21_147 ();
 FILLCELL_X1 FILLER_0_21_149 ();
 FILLCELL_X8 FILLER_0_21_155 ();
 FILLCELL_X8 FILLER_0_21_165 ();
 FILLCELL_X4 FILLER_0_21_173 ();
 FILLCELL_X2 FILLER_0_21_177 ();
 FILLCELL_X1 FILLER_0_21_179 ();
 FILLCELL_X32 FILLER_0_21_201 ();
 FILLCELL_X4 FILLER_0_21_233 ();
 FILLCELL_X2 FILLER_0_21_237 ();
 FILLCELL_X4 FILLER_0_21_241 ();
 FILLCELL_X4 FILLER_0_21_248 ();
 FILLCELL_X2 FILLER_0_21_252 ();
 FILLCELL_X4 FILLER_0_21_257 ();
 FILLCELL_X1 FILLER_0_21_263 ();
 FILLCELL_X2 FILLER_0_21_273 ();
 FILLCELL_X1 FILLER_0_21_297 ();
 FILLCELL_X8 FILLER_0_21_303 ();
 FILLCELL_X2 FILLER_0_21_311 ();
 FILLCELL_X1 FILLER_0_21_318 ();
 FILLCELL_X2 FILLER_0_21_339 ();
 FILLCELL_X2 FILLER_0_21_387 ();
 FILLCELL_X4 FILLER_0_22_1 ();
 FILLCELL_X1 FILLER_0_22_5 ();
 FILLCELL_X8 FILLER_0_22_9 ();
 FILLCELL_X1 FILLER_0_22_17 ();
 FILLCELL_X4 FILLER_0_22_24 ();
 FILLCELL_X1 FILLER_0_22_28 ();
 FILLCELL_X32 FILLER_0_22_32 ();
 FILLCELL_X2 FILLER_0_22_70 ();
 FILLCELL_X2 FILLER_0_22_83 ();
 FILLCELL_X4 FILLER_0_22_98 ();
 FILLCELL_X8 FILLER_0_22_108 ();
 FILLCELL_X1 FILLER_0_22_116 ();
 FILLCELL_X8 FILLER_0_22_125 ();
 FILLCELL_X2 FILLER_0_22_133 ();
 FILLCELL_X1 FILLER_0_22_138 ();
 FILLCELL_X2 FILLER_0_22_144 ();
 FILLCELL_X1 FILLER_0_22_146 ();
 FILLCELL_X2 FILLER_0_22_157 ();
 FILLCELL_X2 FILLER_0_22_171 ();
 FILLCELL_X4 FILLER_0_22_186 ();
 FILLCELL_X2 FILLER_0_22_190 ();
 FILLCELL_X8 FILLER_0_22_218 ();
 FILLCELL_X1 FILLER_0_22_226 ();
 FILLCELL_X2 FILLER_0_22_243 ();
 FILLCELL_X1 FILLER_0_22_245 ();
 FILLCELL_X4 FILLER_0_22_249 ();
 FILLCELL_X2 FILLER_0_22_253 ();
 FILLCELL_X2 FILLER_0_22_286 ();
 FILLCELL_X2 FILLER_0_22_297 ();
 FILLCELL_X1 FILLER_0_22_299 ();
 FILLCELL_X8 FILLER_0_22_305 ();
 FILLCELL_X4 FILLER_0_22_313 ();
 FILLCELL_X1 FILLER_0_22_317 ();
 FILLCELL_X8 FILLER_0_22_323 ();
 FILLCELL_X2 FILLER_0_22_331 ();
 FILLCELL_X2 FILLER_0_22_345 ();
 FILLCELL_X2 FILLER_0_22_381 ();
 FILLCELL_X1 FILLER_0_22_383 ();
 FILLCELL_X1 FILLER_0_23_1 ();
 FILLCELL_X2 FILLER_0_23_10 ();
 FILLCELL_X1 FILLER_0_23_12 ();
 FILLCELL_X1 FILLER_0_23_16 ();
 FILLCELL_X2 FILLER_0_23_19 ();
 FILLCELL_X8 FILLER_0_23_24 ();
 FILLCELL_X2 FILLER_0_23_32 ();
 FILLCELL_X1 FILLER_0_23_34 ();
 FILLCELL_X1 FILLER_0_23_45 ();
 FILLCELL_X2 FILLER_0_23_49 ();
 FILLCELL_X1 FILLER_0_23_51 ();
 FILLCELL_X2 FILLER_0_23_58 ();
 FILLCELL_X1 FILLER_0_23_78 ();
 FILLCELL_X2 FILLER_0_23_85 ();
 FILLCELL_X1 FILLER_0_23_87 ();
 FILLCELL_X4 FILLER_0_23_91 ();
 FILLCELL_X1 FILLER_0_23_95 ();
 FILLCELL_X8 FILLER_0_23_98 ();
 FILLCELL_X2 FILLER_0_23_106 ();
 FILLCELL_X1 FILLER_0_23_108 ();
 FILLCELL_X8 FILLER_0_23_115 ();
 FILLCELL_X1 FILLER_0_23_123 ();
 FILLCELL_X8 FILLER_0_23_126 ();
 FILLCELL_X4 FILLER_0_23_134 ();
 FILLCELL_X1 FILLER_0_23_140 ();
 FILLCELL_X1 FILLER_0_23_147 ();
 FILLCELL_X1 FILLER_0_23_170 ();
 FILLCELL_X1 FILLER_0_23_174 ();
 FILLCELL_X16 FILLER_0_23_184 ();
 FILLCELL_X4 FILLER_0_23_200 ();
 FILLCELL_X2 FILLER_0_23_204 ();
 FILLCELL_X1 FILLER_0_23_206 ();
 FILLCELL_X1 FILLER_0_23_210 ();
 FILLCELL_X1 FILLER_0_23_214 ();
 FILLCELL_X1 FILLER_0_23_220 ();
 FILLCELL_X2 FILLER_0_23_223 ();
 FILLCELL_X1 FILLER_0_23_225 ();
 FILLCELL_X2 FILLER_0_23_228 ();
 FILLCELL_X2 FILLER_0_23_233 ();
 FILLCELL_X1 FILLER_0_23_235 ();
 FILLCELL_X2 FILLER_0_23_239 ();
 FILLCELL_X4 FILLER_0_23_249 ();
 FILLCELL_X1 FILLER_0_23_253 ();
 FILLCELL_X2 FILLER_0_23_257 ();
 FILLCELL_X1 FILLER_0_23_284 ();
 FILLCELL_X8 FILLER_0_23_298 ();
 FILLCELL_X4 FILLER_0_23_306 ();
 FILLCELL_X1 FILLER_0_23_310 ();
 FILLCELL_X1 FILLER_0_23_329 ();
 FILLCELL_X1 FILLER_0_23_366 ();
 FILLCELL_X1 FILLER_0_23_379 ();
 FILLCELL_X4 FILLER_0_23_387 ();
 FILLCELL_X1 FILLER_0_23_391 ();
 FILLCELL_X4 FILLER_0_23_397 ();
 FILLCELL_X1 FILLER_0_23_401 ();
 FILLCELL_X4 FILLER_0_23_404 ();
 FILLCELL_X2 FILLER_0_24_1 ();
 FILLCELL_X1 FILLER_0_24_3 ();
 FILLCELL_X2 FILLER_0_24_10 ();
 FILLCELL_X1 FILLER_0_24_12 ();
 FILLCELL_X1 FILLER_0_24_19 ();
 FILLCELL_X2 FILLER_0_24_23 ();
 FILLCELL_X1 FILLER_0_24_25 ();
 FILLCELL_X1 FILLER_0_24_29 ();
 FILLCELL_X8 FILLER_0_24_36 ();
 FILLCELL_X1 FILLER_0_24_44 ();
 FILLCELL_X8 FILLER_0_24_48 ();
 FILLCELL_X4 FILLER_0_24_56 ();
 FILLCELL_X1 FILLER_0_24_60 ();
 FILLCELL_X8 FILLER_0_24_66 ();
 FILLCELL_X2 FILLER_0_24_74 ();
 FILLCELL_X2 FILLER_0_24_78 ();
 FILLCELL_X1 FILLER_0_24_80 ();
 FILLCELL_X2 FILLER_0_24_103 ();
 FILLCELL_X1 FILLER_0_24_105 ();
 FILLCELL_X1 FILLER_0_24_108 ();
 FILLCELL_X1 FILLER_0_24_156 ();
 FILLCELL_X2 FILLER_0_24_163 ();
 FILLCELL_X1 FILLER_0_24_165 ();
 FILLCELL_X2 FILLER_0_24_168 ();
 FILLCELL_X1 FILLER_0_24_170 ();
 FILLCELL_X4 FILLER_0_24_177 ();
 FILLCELL_X16 FILLER_0_24_188 ();
 FILLCELL_X4 FILLER_0_24_204 ();
 FILLCELL_X1 FILLER_0_24_208 ();
 FILLCELL_X4 FILLER_0_24_211 ();
 FILLCELL_X1 FILLER_0_24_225 ();
 FILLCELL_X2 FILLER_0_24_235 ();
 FILLCELL_X1 FILLER_0_24_245 ();
 FILLCELL_X2 FILLER_0_24_253 ();
 FILLCELL_X1 FILLER_0_24_255 ();
 FILLCELL_X2 FILLER_0_24_264 ();
 FILLCELL_X1 FILLER_0_24_266 ();
 FILLCELL_X32 FILLER_0_24_285 ();
 FILLCELL_X4 FILLER_0_24_317 ();
 FILLCELL_X1 FILLER_0_24_336 ();
 FILLCELL_X1 FILLER_0_24_373 ();
 FILLCELL_X2 FILLER_0_24_396 ();
 FILLCELL_X4 FILLER_0_24_400 ();
 FILLCELL_X1 FILLER_0_24_404 ();
 FILLCELL_X2 FILLER_0_25_6 ();
 FILLCELL_X1 FILLER_0_25_8 ();
 FILLCELL_X8 FILLER_0_25_14 ();
 FILLCELL_X4 FILLER_0_25_22 ();
 FILLCELL_X2 FILLER_0_25_26 ();
 FILLCELL_X2 FILLER_0_25_31 ();
 FILLCELL_X1 FILLER_0_25_33 ();
 FILLCELL_X1 FILLER_0_25_63 ();
 FILLCELL_X4 FILLER_0_25_74 ();
 FILLCELL_X2 FILLER_0_25_78 ();
 FILLCELL_X1 FILLER_0_25_80 ();
 FILLCELL_X4 FILLER_0_25_83 ();
 FILLCELL_X2 FILLER_0_25_87 ();
 FILLCELL_X4 FILLER_0_25_104 ();
 FILLCELL_X4 FILLER_0_25_160 ();
 FILLCELL_X2 FILLER_0_25_164 ();
 FILLCELL_X8 FILLER_0_25_189 ();
 FILLCELL_X2 FILLER_0_25_197 ();
 FILLCELL_X1 FILLER_0_25_201 ();
 FILLCELL_X1 FILLER_0_25_204 ();
 FILLCELL_X1 FILLER_0_25_209 ();
 FILLCELL_X1 FILLER_0_25_213 ();
 FILLCELL_X8 FILLER_0_25_217 ();
 FILLCELL_X2 FILLER_0_25_225 ();
 FILLCELL_X1 FILLER_0_25_227 ();
 FILLCELL_X2 FILLER_0_25_234 ();
 FILLCELL_X1 FILLER_0_25_236 ();
 FILLCELL_X2 FILLER_0_25_250 ();
 FILLCELL_X2 FILLER_0_25_260 ();
 FILLCELL_X1 FILLER_0_25_266 ();
 FILLCELL_X2 FILLER_0_25_308 ();
 FILLCELL_X1 FILLER_0_25_310 ();
 FILLCELL_X4 FILLER_0_25_317 ();
 FILLCELL_X2 FILLER_0_25_321 ();
 FILLCELL_X1 FILLER_0_25_323 ();
 FILLCELL_X1 FILLER_0_25_329 ();
 FILLCELL_X1 FILLER_0_25_332 ();
 FILLCELL_X1 FILLER_0_25_343 ();
 FILLCELL_X1 FILLER_0_25_356 ();
 FILLCELL_X4 FILLER_0_25_366 ();
 FILLCELL_X2 FILLER_0_25_370 ();
 FILLCELL_X1 FILLER_0_25_372 ();
 FILLCELL_X2 FILLER_0_25_389 ();
 FILLCELL_X1 FILLER_0_25_407 ();
 FILLCELL_X2 FILLER_0_26_7 ();
 FILLCELL_X1 FILLER_0_26_13 ();
 FILLCELL_X1 FILLER_0_26_20 ();
 FILLCELL_X1 FILLER_0_26_26 ();
 FILLCELL_X8 FILLER_0_26_52 ();
 FILLCELL_X2 FILLER_0_26_60 ();
 FILLCELL_X2 FILLER_0_26_64 ();
 FILLCELL_X2 FILLER_0_26_74 ();
 FILLCELL_X4 FILLER_0_26_88 ();
 FILLCELL_X1 FILLER_0_26_92 ();
 FILLCELL_X1 FILLER_0_26_95 ();
 FILLCELL_X4 FILLER_0_26_101 ();
 FILLCELL_X1 FILLER_0_26_114 ();
 FILLCELL_X4 FILLER_0_26_123 ();
 FILLCELL_X2 FILLER_0_26_127 ();
 FILLCELL_X1 FILLER_0_26_129 ();
 FILLCELL_X8 FILLER_0_26_171 ();
 FILLCELL_X4 FILLER_0_26_179 ();
 FILLCELL_X1 FILLER_0_26_183 ();
 FILLCELL_X1 FILLER_0_26_208 ();
 FILLCELL_X8 FILLER_0_26_220 ();
 FILLCELL_X2 FILLER_0_26_250 ();
 FILLCELL_X4 FILLER_0_26_258 ();
 FILLCELL_X1 FILLER_0_26_262 ();
 FILLCELL_X1 FILLER_0_26_298 ();
 FILLCELL_X8 FILLER_0_26_322 ();
 FILLCELL_X1 FILLER_0_26_330 ();
 FILLCELL_X8 FILLER_0_26_334 ();
 FILLCELL_X16 FILLER_0_26_370 ();
 FILLCELL_X8 FILLER_0_26_386 ();
 FILLCELL_X8 FILLER_0_26_397 ();
 FILLCELL_X1 FILLER_0_26_405 ();
 FILLCELL_X4 FILLER_0_27_1 ();
 FILLCELL_X1 FILLER_0_27_5 ();
 FILLCELL_X1 FILLER_0_27_9 ();
 FILLCELL_X8 FILLER_0_27_12 ();
 FILLCELL_X4 FILLER_0_27_20 ();
 FILLCELL_X2 FILLER_0_27_24 ();
 FILLCELL_X1 FILLER_0_27_26 ();
 FILLCELL_X2 FILLER_0_27_49 ();
 FILLCELL_X1 FILLER_0_27_51 ();
 FILLCELL_X1 FILLER_0_27_86 ();
 FILLCELL_X2 FILLER_0_27_92 ();
 FILLCELL_X1 FILLER_0_27_96 ();
 FILLCELL_X8 FILLER_0_27_123 ();
 FILLCELL_X4 FILLER_0_27_131 ();
 FILLCELL_X1 FILLER_0_27_135 ();
 FILLCELL_X16 FILLER_0_27_151 ();
 FILLCELL_X4 FILLER_0_27_167 ();
 FILLCELL_X1 FILLER_0_27_171 ();
 FILLCELL_X4 FILLER_0_27_175 ();
 FILLCELL_X2 FILLER_0_27_179 ();
 FILLCELL_X1 FILLER_0_27_181 ();
 FILLCELL_X1 FILLER_0_27_184 ();
 FILLCELL_X2 FILLER_0_27_200 ();
 FILLCELL_X2 FILLER_0_27_221 ();
 FILLCELL_X1 FILLER_0_27_223 ();
 FILLCELL_X1 FILLER_0_27_227 ();
 FILLCELL_X2 FILLER_0_27_231 ();
 FILLCELL_X8 FILLER_0_27_243 ();
 FILLCELL_X4 FILLER_0_27_251 ();
 FILLCELL_X2 FILLER_0_27_257 ();
 FILLCELL_X8 FILLER_0_27_272 ();
 FILLCELL_X1 FILLER_0_27_291 ();
 FILLCELL_X8 FILLER_0_27_294 ();
 FILLCELL_X4 FILLER_0_27_302 ();
 FILLCELL_X1 FILLER_0_27_306 ();
 FILLCELL_X2 FILLER_0_27_331 ();
 FILLCELL_X32 FILLER_0_27_368 ();
 FILLCELL_X8 FILLER_0_27_400 ();
 FILLCELL_X32 FILLER_0_28_1 ();
 FILLCELL_X2 FILLER_0_28_49 ();
 FILLCELL_X1 FILLER_0_28_51 ();
 FILLCELL_X1 FILLER_0_28_68 ();
 FILLCELL_X1 FILLER_0_28_71 ();
 FILLCELL_X1 FILLER_0_28_76 ();
 FILLCELL_X8 FILLER_0_28_80 ();
 FILLCELL_X4 FILLER_0_28_88 ();
 FILLCELL_X2 FILLER_0_28_92 ();
 FILLCELL_X1 FILLER_0_28_94 ();
 FILLCELL_X8 FILLER_0_28_110 ();
 FILLCELL_X4 FILLER_0_28_120 ();
 FILLCELL_X2 FILLER_0_28_124 ();
 FILLCELL_X32 FILLER_0_28_130 ();
 FILLCELL_X4 FILLER_0_28_165 ();
 FILLCELL_X2 FILLER_0_28_169 ();
 FILLCELL_X1 FILLER_0_28_171 ();
 FILLCELL_X1 FILLER_0_28_175 ();
 FILLCELL_X2 FILLER_0_28_181 ();
 FILLCELL_X2 FILLER_0_28_193 ();
 FILLCELL_X4 FILLER_0_28_200 ();
 FILLCELL_X1 FILLER_0_28_206 ();
 FILLCELL_X8 FILLER_0_28_211 ();
 FILLCELL_X4 FILLER_0_28_219 ();
 FILLCELL_X8 FILLER_0_28_236 ();
 FILLCELL_X2 FILLER_0_28_244 ();
 FILLCELL_X1 FILLER_0_28_246 ();
 FILLCELL_X4 FILLER_0_28_250 ();
 FILLCELL_X1 FILLER_0_28_257 ();
 FILLCELL_X2 FILLER_0_28_271 ();
 FILLCELL_X1 FILLER_0_28_273 ();
 FILLCELL_X4 FILLER_0_28_280 ();
 FILLCELL_X2 FILLER_0_28_284 ();
 FILLCELL_X1 FILLER_0_28_286 ();
 FILLCELL_X8 FILLER_0_28_296 ();
 FILLCELL_X4 FILLER_0_28_304 ();
 FILLCELL_X2 FILLER_0_28_308 ();
 FILLCELL_X4 FILLER_0_28_317 ();
 FILLCELL_X4 FILLER_0_28_324 ();
 FILLCELL_X1 FILLER_0_28_328 ();
 FILLCELL_X4 FILLER_0_28_331 ();
 FILLCELL_X2 FILLER_0_28_335 ();
 FILLCELL_X1 FILLER_0_28_337 ();
 FILLCELL_X2 FILLER_0_28_355 ();
 FILLCELL_X16 FILLER_0_28_359 ();
 FILLCELL_X4 FILLER_0_28_375 ();
 FILLCELL_X1 FILLER_0_28_379 ();
 FILLCELL_X16 FILLER_0_28_389 ();
 FILLCELL_X2 FILLER_0_28_405 ();
 FILLCELL_X1 FILLER_0_28_407 ();
 FILLCELL_X32 FILLER_0_29_1 ();
 FILLCELL_X2 FILLER_0_29_33 ();
 FILLCELL_X1 FILLER_0_29_35 ();
 FILLCELL_X8 FILLER_0_29_46 ();
 FILLCELL_X4 FILLER_0_29_54 ();
 FILLCELL_X1 FILLER_0_29_69 ();
 FILLCELL_X1 FILLER_0_29_90 ();
 FILLCELL_X1 FILLER_0_29_132 ();
 FILLCELL_X2 FILLER_0_29_138 ();
 FILLCELL_X1 FILLER_0_29_140 ();
 FILLCELL_X8 FILLER_0_29_149 ();
 FILLCELL_X4 FILLER_0_29_157 ();
 FILLCELL_X1 FILLER_0_29_167 ();
 FILLCELL_X2 FILLER_0_29_177 ();
 FILLCELL_X16 FILLER_0_29_182 ();
 FILLCELL_X1 FILLER_0_29_198 ();
 FILLCELL_X2 FILLER_0_29_235 ();
 FILLCELL_X2 FILLER_0_29_240 ();
 FILLCELL_X1 FILLER_0_29_242 ();
 FILLCELL_X1 FILLER_0_29_258 ();
 FILLCELL_X1 FILLER_0_29_266 ();
 FILLCELL_X4 FILLER_0_29_274 ();
 FILLCELL_X2 FILLER_0_29_278 ();
 FILLCELL_X1 FILLER_0_29_280 ();
 FILLCELL_X2 FILLER_0_29_303 ();
 FILLCELL_X1 FILLER_0_29_309 ();
 FILLCELL_X4 FILLER_0_29_329 ();
 FILLCELL_X1 FILLER_0_29_333 ();
 FILLCELL_X2 FILLER_0_29_341 ();
 FILLCELL_X1 FILLER_0_29_350 ();
 FILLCELL_X1 FILLER_0_29_353 ();
 FILLCELL_X1 FILLER_0_29_357 ();
 FILLCELL_X4 FILLER_0_29_369 ();
 FILLCELL_X2 FILLER_0_29_373 ();
 FILLCELL_X1 FILLER_0_29_375 ();
 FILLCELL_X1 FILLER_0_29_381 ();
 FILLCELL_X8 FILLER_0_29_394 ();
 FILLCELL_X4 FILLER_0_29_402 ();
 FILLCELL_X2 FILLER_0_29_406 ();
 FILLCELL_X32 FILLER_0_30_1 ();
 FILLCELL_X16 FILLER_0_30_33 ();
 FILLCELL_X4 FILLER_0_30_81 ();
 FILLCELL_X1 FILLER_0_30_85 ();
 FILLCELL_X1 FILLER_0_30_102 ();
 FILLCELL_X1 FILLER_0_30_106 ();
 FILLCELL_X1 FILLER_0_30_114 ();
 FILLCELL_X8 FILLER_0_30_144 ();
 FILLCELL_X2 FILLER_0_30_152 ();
 FILLCELL_X1 FILLER_0_30_157 ();
 FILLCELL_X4 FILLER_0_30_166 ();
 FILLCELL_X2 FILLER_0_30_170 ();
 FILLCELL_X16 FILLER_0_30_180 ();
 FILLCELL_X1 FILLER_0_30_196 ();
 FILLCELL_X8 FILLER_0_30_211 ();
 FILLCELL_X4 FILLER_0_30_219 ();
 FILLCELL_X1 FILLER_0_30_223 ();
 FILLCELL_X8 FILLER_0_30_237 ();
 FILLCELL_X4 FILLER_0_30_245 ();
 FILLCELL_X1 FILLER_0_30_255 ();
 FILLCELL_X16 FILLER_0_30_264 ();
 FILLCELL_X2 FILLER_0_30_280 ();
 FILLCELL_X2 FILLER_0_30_289 ();
 FILLCELL_X2 FILLER_0_30_294 ();
 FILLCELL_X1 FILLER_0_30_296 ();
 FILLCELL_X8 FILLER_0_30_305 ();
 FILLCELL_X2 FILLER_0_30_316 ();
 FILLCELL_X1 FILLER_0_30_330 ();
 FILLCELL_X2 FILLER_0_30_336 ();
 FILLCELL_X1 FILLER_0_30_345 ();
 FILLCELL_X4 FILLER_0_30_349 ();
 FILLCELL_X8 FILLER_0_30_369 ();
 FILLCELL_X4 FILLER_0_30_402 ();
 FILLCELL_X2 FILLER_0_30_406 ();
 FILLCELL_X32 FILLER_0_31_1 ();
 FILLCELL_X16 FILLER_0_31_33 ();
 FILLCELL_X8 FILLER_0_31_49 ();
 FILLCELL_X4 FILLER_0_31_57 ();
 FILLCELL_X1 FILLER_0_31_61 ();
 FILLCELL_X1 FILLER_0_31_64 ();
 FILLCELL_X8 FILLER_0_31_78 ();
 FILLCELL_X4 FILLER_0_31_86 ();
 FILLCELL_X2 FILLER_0_31_90 ();
 FILLCELL_X1 FILLER_0_31_92 ();
 FILLCELL_X4 FILLER_0_31_122 ();
 FILLCELL_X2 FILLER_0_31_126 ();
 FILLCELL_X1 FILLER_0_31_128 ();
 FILLCELL_X8 FILLER_0_31_131 ();
 FILLCELL_X4 FILLER_0_31_139 ();
 FILLCELL_X2 FILLER_0_31_143 ();
 FILLCELL_X1 FILLER_0_31_145 ();
 FILLCELL_X4 FILLER_0_31_153 ();
 FILLCELL_X2 FILLER_0_31_170 ();
 FILLCELL_X2 FILLER_0_31_184 ();
 FILLCELL_X1 FILLER_0_31_186 ();
 FILLCELL_X4 FILLER_0_31_190 ();
 FILLCELL_X1 FILLER_0_31_194 ();
 FILLCELL_X1 FILLER_0_31_198 ();
 FILLCELL_X2 FILLER_0_31_212 ();
 FILLCELL_X2 FILLER_0_31_217 ();
 FILLCELL_X1 FILLER_0_31_219 ();
 FILLCELL_X2 FILLER_0_31_225 ();
 FILLCELL_X2 FILLER_0_31_230 ();
 FILLCELL_X4 FILLER_0_31_236 ();
 FILLCELL_X2 FILLER_0_31_240 ();
 FILLCELL_X1 FILLER_0_31_242 ();
 FILLCELL_X2 FILLER_0_31_260 ();
 FILLCELL_X4 FILLER_0_31_272 ();
 FILLCELL_X2 FILLER_0_31_276 ();
 FILLCELL_X1 FILLER_0_31_285 ();
 FILLCELL_X4 FILLER_0_31_292 ();
 FILLCELL_X2 FILLER_0_31_296 ();
 FILLCELL_X1 FILLER_0_31_298 ();
 FILLCELL_X16 FILLER_0_31_302 ();
 FILLCELL_X1 FILLER_0_31_318 ();
 FILLCELL_X2 FILLER_0_31_339 ();
 FILLCELL_X1 FILLER_0_31_341 ();
 FILLCELL_X2 FILLER_0_31_365 ();
 FILLCELL_X2 FILLER_0_31_372 ();
 FILLCELL_X1 FILLER_0_31_374 ();
 FILLCELL_X1 FILLER_0_31_380 ();
 FILLCELL_X2 FILLER_0_31_387 ();
 FILLCELL_X1 FILLER_0_31_389 ();
 FILLCELL_X2 FILLER_0_31_397 ();
 FILLCELL_X1 FILLER_0_31_399 ();
 FILLCELL_X2 FILLER_0_31_403 ();
 FILLCELL_X32 FILLER_0_32_1 ();
 FILLCELL_X32 FILLER_0_32_33 ();
 FILLCELL_X32 FILLER_0_32_65 ();
 FILLCELL_X4 FILLER_0_32_97 ();
 FILLCELL_X2 FILLER_0_32_101 ();
 FILLCELL_X4 FILLER_0_32_105 ();
 FILLCELL_X1 FILLER_0_32_109 ();
 FILLCELL_X32 FILLER_0_32_112 ();
 FILLCELL_X8 FILLER_0_32_144 ();
 FILLCELL_X4 FILLER_0_32_152 ();
 FILLCELL_X2 FILLER_0_32_168 ();
 FILLCELL_X1 FILLER_0_32_170 ();
 FILLCELL_X2 FILLER_0_32_175 ();
 FILLCELL_X1 FILLER_0_32_177 ();
 FILLCELL_X4 FILLER_0_32_181 ();
 FILLCELL_X2 FILLER_0_32_185 ();
 FILLCELL_X2 FILLER_0_32_202 ();
 FILLCELL_X4 FILLER_0_32_208 ();
 FILLCELL_X2 FILLER_0_32_221 ();
 FILLCELL_X1 FILLER_0_32_223 ();
 FILLCELL_X2 FILLER_0_32_229 ();
 FILLCELL_X1 FILLER_0_32_231 ();
 FILLCELL_X2 FILLER_0_32_235 ();
 FILLCELL_X1 FILLER_0_32_237 ();
 FILLCELL_X4 FILLER_0_32_241 ();
 FILLCELL_X1 FILLER_0_32_245 ();
 FILLCELL_X1 FILLER_0_32_249 ();
 FILLCELL_X1 FILLER_0_32_254 ();
 FILLCELL_X2 FILLER_0_32_295 ();
 FILLCELL_X1 FILLER_0_32_301 ();
 FILLCELL_X1 FILLER_0_32_306 ();
 FILLCELL_X1 FILLER_0_32_311 ();
 FILLCELL_X1 FILLER_0_32_316 ();
 FILLCELL_X1 FILLER_0_32_320 ();
 FILLCELL_X4 FILLER_0_32_325 ();
 FILLCELL_X8 FILLER_0_32_332 ();
 FILLCELL_X1 FILLER_0_32_364 ();
 FILLCELL_X4 FILLER_0_32_368 ();
 FILLCELL_X2 FILLER_0_32_372 ();
 FILLCELL_X1 FILLER_0_32_374 ();
 FILLCELL_X1 FILLER_0_32_383 ();
 FILLCELL_X1 FILLER_0_32_404 ();
 FILLCELL_X32 FILLER_0_33_1 ();
 FILLCELL_X32 FILLER_0_33_33 ();
 FILLCELL_X32 FILLER_0_33_65 ();
 FILLCELL_X32 FILLER_0_33_97 ();
 FILLCELL_X16 FILLER_0_33_129 ();
 FILLCELL_X8 FILLER_0_33_145 ();
 FILLCELL_X2 FILLER_0_33_153 ();
 FILLCELL_X1 FILLER_0_33_155 ();
 FILLCELL_X2 FILLER_0_33_173 ();
 FILLCELL_X1 FILLER_0_33_182 ();
 FILLCELL_X1 FILLER_0_33_193 ();
 FILLCELL_X4 FILLER_0_33_207 ();
 FILLCELL_X1 FILLER_0_33_211 ();
 FILLCELL_X1 FILLER_0_33_224 ();
 FILLCELL_X4 FILLER_0_33_228 ();
 FILLCELL_X4 FILLER_0_33_235 ();
 FILLCELL_X2 FILLER_0_33_245 ();
 FILLCELL_X1 FILLER_0_33_247 ();
 FILLCELL_X16 FILLER_0_33_251 ();
 FILLCELL_X2 FILLER_0_33_267 ();
 FILLCELL_X1 FILLER_0_33_269 ();
 FILLCELL_X4 FILLER_0_33_274 ();
 FILLCELL_X2 FILLER_0_33_278 ();
 FILLCELL_X1 FILLER_0_33_280 ();
 FILLCELL_X1 FILLER_0_33_291 ();
 FILLCELL_X2 FILLER_0_33_300 ();
 FILLCELL_X4 FILLER_0_33_310 ();
 FILLCELL_X1 FILLER_0_33_314 ();
 FILLCELL_X2 FILLER_0_33_318 ();
 FILLCELL_X1 FILLER_0_33_324 ();
 FILLCELL_X4 FILLER_0_33_340 ();
 FILLCELL_X16 FILLER_0_33_351 ();
 FILLCELL_X1 FILLER_0_33_367 ();
 FILLCELL_X1 FILLER_0_33_380 ();
 FILLCELL_X4 FILLER_0_33_385 ();
 FILLCELL_X2 FILLER_0_33_389 ();
 FILLCELL_X1 FILLER_0_33_391 ();
 FILLCELL_X2 FILLER_0_33_402 ();
 FILLCELL_X1 FILLER_0_33_404 ();
 FILLCELL_X32 FILLER_0_34_1 ();
 FILLCELL_X32 FILLER_0_34_33 ();
 FILLCELL_X32 FILLER_0_34_65 ();
 FILLCELL_X32 FILLER_0_34_97 ();
 FILLCELL_X16 FILLER_0_34_129 ();
 FILLCELL_X8 FILLER_0_34_145 ();
 FILLCELL_X2 FILLER_0_34_153 ();
 FILLCELL_X1 FILLER_0_34_155 ();
 FILLCELL_X2 FILLER_0_34_163 ();
 FILLCELL_X16 FILLER_0_34_169 ();
 FILLCELL_X4 FILLER_0_34_185 ();
 FILLCELL_X1 FILLER_0_34_189 ();
 FILLCELL_X1 FILLER_0_34_204 ();
 FILLCELL_X2 FILLER_0_34_210 ();
 FILLCELL_X1 FILLER_0_34_212 ();
 FILLCELL_X1 FILLER_0_34_215 ();
 FILLCELL_X1 FILLER_0_34_219 ();
 FILLCELL_X1 FILLER_0_34_242 ();
 FILLCELL_X1 FILLER_0_34_261 ();
 FILLCELL_X1 FILLER_0_34_265 ();
 FILLCELL_X1 FILLER_0_34_268 ();
 FILLCELL_X4 FILLER_0_34_277 ();
 FILLCELL_X2 FILLER_0_34_281 ();
 FILLCELL_X2 FILLER_0_34_296 ();
 FILLCELL_X1 FILLER_0_34_298 ();
 FILLCELL_X4 FILLER_0_34_315 ();
 FILLCELL_X4 FILLER_0_34_322 ();
 FILLCELL_X2 FILLER_0_34_326 ();
 FILLCELL_X4 FILLER_0_34_331 ();
 FILLCELL_X1 FILLER_0_34_345 ();
 FILLCELL_X1 FILLER_0_34_349 ();
 FILLCELL_X1 FILLER_0_34_354 ();
 FILLCELL_X2 FILLER_0_34_362 ();
 FILLCELL_X1 FILLER_0_34_364 ();
 FILLCELL_X1 FILLER_0_34_388 ();
 FILLCELL_X2 FILLER_0_34_406 ();
 FILLCELL_X32 FILLER_0_35_1 ();
 FILLCELL_X32 FILLER_0_35_33 ();
 FILLCELL_X32 FILLER_0_35_65 ();
 FILLCELL_X32 FILLER_0_35_97 ();
 FILLCELL_X16 FILLER_0_35_129 ();
 FILLCELL_X8 FILLER_0_35_145 ();
 FILLCELL_X8 FILLER_0_35_166 ();
 FILLCELL_X4 FILLER_0_35_174 ();
 FILLCELL_X2 FILLER_0_35_178 ();
 FILLCELL_X2 FILLER_0_35_192 ();
 FILLCELL_X1 FILLER_0_35_194 ();
 FILLCELL_X4 FILLER_0_35_202 ();
 FILLCELL_X2 FILLER_0_35_206 ();
 FILLCELL_X1 FILLER_0_35_208 ();
 FILLCELL_X1 FILLER_0_35_214 ();
 FILLCELL_X8 FILLER_0_35_218 ();
 FILLCELL_X2 FILLER_0_35_226 ();
 FILLCELL_X1 FILLER_0_35_233 ();
 FILLCELL_X1 FILLER_0_35_241 ();
 FILLCELL_X4 FILLER_0_35_250 ();
 FILLCELL_X2 FILLER_0_35_254 ();
 FILLCELL_X1 FILLER_0_35_256 ();
 FILLCELL_X1 FILLER_0_35_260 ();
 FILLCELL_X4 FILLER_0_35_264 ();
 FILLCELL_X2 FILLER_0_35_268 ();
 FILLCELL_X4 FILLER_0_35_282 ();
 FILLCELL_X4 FILLER_0_35_293 ();
 FILLCELL_X2 FILLER_0_35_297 ();
 FILLCELL_X1 FILLER_0_35_299 ();
 FILLCELL_X2 FILLER_0_35_305 ();
 FILLCELL_X1 FILLER_0_35_307 ();
 FILLCELL_X4 FILLER_0_35_319 ();
 FILLCELL_X2 FILLER_0_35_323 ();
 FILLCELL_X4 FILLER_0_35_329 ();
 FILLCELL_X2 FILLER_0_35_349 ();
 FILLCELL_X2 FILLER_0_35_355 ();
 FILLCELL_X8 FILLER_0_35_360 ();
 FILLCELL_X2 FILLER_0_35_368 ();
 FILLCELL_X16 FILLER_0_35_379 ();
 FILLCELL_X1 FILLER_0_35_402 ();
 FILLCELL_X2 FILLER_0_35_406 ();
 FILLCELL_X32 FILLER_0_36_1 ();
 FILLCELL_X32 FILLER_0_36_33 ();
 FILLCELL_X32 FILLER_0_36_65 ();
 FILLCELL_X32 FILLER_0_36_97 ();
 FILLCELL_X16 FILLER_0_36_129 ();
 FILLCELL_X4 FILLER_0_36_145 ();
 FILLCELL_X1 FILLER_0_36_159 ();
 FILLCELL_X2 FILLER_0_36_163 ();
 FILLCELL_X1 FILLER_0_36_168 ();
 FILLCELL_X2 FILLER_0_36_173 ();
 FILLCELL_X2 FILLER_0_36_181 ();
 FILLCELL_X1 FILLER_0_36_186 ();
 FILLCELL_X8 FILLER_0_36_191 ();
 FILLCELL_X4 FILLER_0_36_199 ();
 FILLCELL_X1 FILLER_0_36_223 ();
 FILLCELL_X4 FILLER_0_36_226 ();
 FILLCELL_X2 FILLER_0_36_230 ();
 FILLCELL_X1 FILLER_0_36_232 ();
 FILLCELL_X8 FILLER_0_36_235 ();
 FILLCELL_X2 FILLER_0_36_243 ();
 FILLCELL_X2 FILLER_0_36_257 ();
 FILLCELL_X4 FILLER_0_36_262 ();
 FILLCELL_X1 FILLER_0_36_266 ();
 FILLCELL_X8 FILLER_0_36_282 ();
 FILLCELL_X1 FILLER_0_36_290 ();
 FILLCELL_X1 FILLER_0_36_299 ();
 FILLCELL_X8 FILLER_0_36_311 ();
 FILLCELL_X2 FILLER_0_36_319 ();
 FILLCELL_X1 FILLER_0_36_348 ();
 FILLCELL_X1 FILLER_0_36_355 ();
 FILLCELL_X8 FILLER_0_36_359 ();
 FILLCELL_X4 FILLER_0_36_367 ();
 FILLCELL_X8 FILLER_0_36_382 ();
 FILLCELL_X2 FILLER_0_36_390 ();
 FILLCELL_X1 FILLER_0_36_392 ();
 FILLCELL_X32 FILLER_0_37_1 ();
 FILLCELL_X32 FILLER_0_37_33 ();
 FILLCELL_X32 FILLER_0_37_65 ();
 FILLCELL_X32 FILLER_0_37_97 ();
 FILLCELL_X16 FILLER_0_37_129 ();
 FILLCELL_X8 FILLER_0_37_145 ();
 FILLCELL_X4 FILLER_0_37_153 ();
 FILLCELL_X2 FILLER_0_37_157 ();
 FILLCELL_X1 FILLER_0_37_159 ();
 FILLCELL_X4 FILLER_0_37_182 ();
 FILLCELL_X1 FILLER_0_37_186 ();
 FILLCELL_X4 FILLER_0_37_194 ();
 FILLCELL_X1 FILLER_0_37_198 ();
 FILLCELL_X1 FILLER_0_37_212 ();
 FILLCELL_X2 FILLER_0_37_216 ();
 FILLCELL_X4 FILLER_0_37_221 ();
 FILLCELL_X2 FILLER_0_37_225 ();
 FILLCELL_X2 FILLER_0_37_240 ();
 FILLCELL_X1 FILLER_0_37_244 ();
 FILLCELL_X1 FILLER_0_37_248 ();
 FILLCELL_X2 FILLER_0_37_253 ();
 FILLCELL_X2 FILLER_0_37_262 ();
 FILLCELL_X1 FILLER_0_37_264 ();
 FILLCELL_X16 FILLER_0_37_275 ();
 FILLCELL_X4 FILLER_0_37_291 ();
 FILLCELL_X2 FILLER_0_37_295 ();
 FILLCELL_X2 FILLER_0_37_302 ();
 FILLCELL_X1 FILLER_0_37_304 ();
 FILLCELL_X2 FILLER_0_37_314 ();
 FILLCELL_X1 FILLER_0_37_316 ();
 FILLCELL_X2 FILLER_0_37_319 ();
 FILLCELL_X2 FILLER_0_37_324 ();
 FILLCELL_X1 FILLER_0_37_326 ();
 FILLCELL_X4 FILLER_0_37_365 ();
 FILLCELL_X2 FILLER_0_37_390 ();
 FILLCELL_X2 FILLER_0_37_406 ();
 FILLCELL_X32 FILLER_0_38_1 ();
 FILLCELL_X32 FILLER_0_38_33 ();
 FILLCELL_X32 FILLER_0_38_65 ();
 FILLCELL_X32 FILLER_0_38_97 ();
 FILLCELL_X32 FILLER_0_38_129 ();
 FILLCELL_X1 FILLER_0_38_161 ();
 FILLCELL_X2 FILLER_0_38_172 ();
 FILLCELL_X2 FILLER_0_38_182 ();
 FILLCELL_X8 FILLER_0_38_195 ();
 FILLCELL_X4 FILLER_0_38_203 ();
 FILLCELL_X2 FILLER_0_38_207 ();
 FILLCELL_X1 FILLER_0_38_218 ();
 FILLCELL_X8 FILLER_0_38_222 ();
 FILLCELL_X1 FILLER_0_38_230 ();
 FILLCELL_X2 FILLER_0_38_234 ();
 FILLCELL_X4 FILLER_0_38_242 ();
 FILLCELL_X8 FILLER_0_38_249 ();
 FILLCELL_X1 FILLER_0_38_257 ();
 FILLCELL_X8 FILLER_0_38_260 ();
 FILLCELL_X4 FILLER_0_38_286 ();
 FILLCELL_X2 FILLER_0_38_290 ();
 FILLCELL_X1 FILLER_0_38_292 ();
 FILLCELL_X8 FILLER_0_38_297 ();
 FILLCELL_X2 FILLER_0_38_305 ();
 FILLCELL_X1 FILLER_0_38_307 ();
 FILLCELL_X16 FILLER_0_38_324 ();
 FILLCELL_X2 FILLER_0_38_340 ();
 FILLCELL_X8 FILLER_0_38_365 ();
 FILLCELL_X2 FILLER_0_38_373 ();
 FILLCELL_X16 FILLER_0_38_377 ();
 FILLCELL_X2 FILLER_0_38_393 ();
 FILLCELL_X1 FILLER_0_38_395 ();
 FILLCELL_X32 FILLER_0_39_1 ();
 FILLCELL_X32 FILLER_0_39_33 ();
 FILLCELL_X32 FILLER_0_39_65 ();
 FILLCELL_X32 FILLER_0_39_97 ();
 FILLCELL_X32 FILLER_0_39_129 ();
 FILLCELL_X32 FILLER_0_39_161 ();
 FILLCELL_X16 FILLER_0_39_193 ();
 FILLCELL_X4 FILLER_0_39_209 ();
 FILLCELL_X2 FILLER_0_39_213 ();
 FILLCELL_X2 FILLER_0_39_218 ();
 FILLCELL_X8 FILLER_0_39_222 ();
 FILLCELL_X2 FILLER_0_39_230 ();
 FILLCELL_X4 FILLER_0_39_244 ();
 FILLCELL_X2 FILLER_0_39_262 ();
 FILLCELL_X1 FILLER_0_39_264 ();
 FILLCELL_X2 FILLER_0_39_268 ();
 FILLCELL_X1 FILLER_0_39_270 ();
 FILLCELL_X1 FILLER_0_39_278 ();
 FILLCELL_X8 FILLER_0_39_283 ();
 FILLCELL_X1 FILLER_0_39_291 ();
 FILLCELL_X4 FILLER_0_39_306 ();
 FILLCELL_X2 FILLER_0_39_310 ();
 FILLCELL_X8 FILLER_0_39_322 ();
 FILLCELL_X1 FILLER_0_39_330 ();
 FILLCELL_X2 FILLER_0_39_338 ();
 FILLCELL_X4 FILLER_0_39_364 ();
 FILLCELL_X1 FILLER_0_39_404 ();
 FILLCELL_X32 FILLER_0_40_1 ();
 FILLCELL_X32 FILLER_0_40_33 ();
 FILLCELL_X32 FILLER_0_40_65 ();
 FILLCELL_X32 FILLER_0_40_97 ();
 FILLCELL_X32 FILLER_0_40_129 ();
 FILLCELL_X32 FILLER_0_40_161 ();
 FILLCELL_X16 FILLER_0_40_193 ();
 FILLCELL_X2 FILLER_0_40_209 ();
 FILLCELL_X1 FILLER_0_40_211 ();
 FILLCELL_X8 FILLER_0_40_222 ();
 FILLCELL_X1 FILLER_0_40_230 ();
 FILLCELL_X2 FILLER_0_40_239 ();
 FILLCELL_X1 FILLER_0_40_241 ();
 FILLCELL_X1 FILLER_0_40_250 ();
 FILLCELL_X1 FILLER_0_40_286 ();
 FILLCELL_X1 FILLER_0_40_305 ();
 FILLCELL_X2 FILLER_0_40_313 ();
 FILLCELL_X2 FILLER_0_40_319 ();
 FILLCELL_X1 FILLER_0_40_321 ();
 FILLCELL_X8 FILLER_0_40_325 ();
 FILLCELL_X2 FILLER_0_40_333 ();
 FILLCELL_X1 FILLER_0_40_335 ();
 FILLCELL_X1 FILLER_0_40_338 ();
 FILLCELL_X1 FILLER_0_40_355 ();
 FILLCELL_X8 FILLER_0_40_359 ();
 FILLCELL_X8 FILLER_0_40_379 ();
 FILLCELL_X4 FILLER_0_40_387 ();
 FILLCELL_X1 FILLER_0_40_391 ();
 FILLCELL_X2 FILLER_0_40_405 ();
 FILLCELL_X1 FILLER_0_40_407 ();
 FILLCELL_X32 FILLER_0_41_1 ();
 FILLCELL_X32 FILLER_0_41_33 ();
 FILLCELL_X32 FILLER_0_41_65 ();
 FILLCELL_X32 FILLER_0_41_97 ();
 FILLCELL_X32 FILLER_0_41_129 ();
 FILLCELL_X32 FILLER_0_41_161 ();
 FILLCELL_X1 FILLER_0_41_193 ();
 FILLCELL_X8 FILLER_0_41_203 ();
 FILLCELL_X2 FILLER_0_41_211 ();
 FILLCELL_X1 FILLER_0_41_213 ();
 FILLCELL_X2 FILLER_0_41_233 ();
 FILLCELL_X8 FILLER_0_41_246 ();
 FILLCELL_X4 FILLER_0_41_262 ();
 FILLCELL_X1 FILLER_0_41_266 ();
 FILLCELL_X8 FILLER_0_41_276 ();
 FILLCELL_X2 FILLER_0_41_284 ();
 FILLCELL_X1 FILLER_0_41_286 ();
 FILLCELL_X2 FILLER_0_41_293 ();
 FILLCELL_X1 FILLER_0_41_298 ();
 FILLCELL_X1 FILLER_0_41_316 ();
 FILLCELL_X2 FILLER_0_41_320 ();
 FILLCELL_X1 FILLER_0_41_334 ();
 FILLCELL_X16 FILLER_0_41_350 ();
 FILLCELL_X8 FILLER_0_41_366 ();
 FILLCELL_X4 FILLER_0_41_390 ();
 FILLCELL_X1 FILLER_0_41_394 ();
 FILLCELL_X32 FILLER_0_42_1 ();
 FILLCELL_X32 FILLER_0_42_33 ();
 FILLCELL_X32 FILLER_0_42_65 ();
 FILLCELL_X32 FILLER_0_42_97 ();
 FILLCELL_X32 FILLER_0_42_129 ();
 FILLCELL_X32 FILLER_0_42_161 ();
 FILLCELL_X8 FILLER_0_42_193 ();
 FILLCELL_X4 FILLER_0_42_201 ();
 FILLCELL_X2 FILLER_0_42_205 ();
 FILLCELL_X1 FILLER_0_42_207 ();
 FILLCELL_X1 FILLER_0_42_265 ();
 FILLCELL_X1 FILLER_0_42_277 ();
 FILLCELL_X1 FILLER_0_42_288 ();
 FILLCELL_X2 FILLER_0_42_299 ();
 FILLCELL_X1 FILLER_0_42_301 ();
 FILLCELL_X8 FILLER_0_42_306 ();
 FILLCELL_X2 FILLER_0_42_317 ();
 FILLCELL_X1 FILLER_0_42_319 ();
 FILLCELL_X4 FILLER_0_42_328 ();
 FILLCELL_X2 FILLER_0_42_332 ();
 FILLCELL_X8 FILLER_0_42_357 ();
 FILLCELL_X1 FILLER_0_42_365 ();
 FILLCELL_X4 FILLER_0_42_370 ();
 FILLCELL_X2 FILLER_0_42_374 ();
 FILLCELL_X16 FILLER_0_42_378 ();
 FILLCELL_X1 FILLER_0_42_394 ();
 FILLCELL_X32 FILLER_0_43_1 ();
 FILLCELL_X32 FILLER_0_43_33 ();
 FILLCELL_X32 FILLER_0_43_65 ();
 FILLCELL_X32 FILLER_0_43_97 ();
 FILLCELL_X32 FILLER_0_43_129 ();
 FILLCELL_X32 FILLER_0_43_161 ();
 FILLCELL_X32 FILLER_0_43_193 ();
 FILLCELL_X4 FILLER_0_43_225 ();
 FILLCELL_X8 FILLER_0_43_233 ();
 FILLCELL_X1 FILLER_0_43_241 ();
 FILLCELL_X1 FILLER_0_43_254 ();
 FILLCELL_X1 FILLER_0_43_259 ();
 FILLCELL_X4 FILLER_0_43_264 ();
 FILLCELL_X2 FILLER_0_43_268 ();
 FILLCELL_X1 FILLER_0_43_270 ();
 FILLCELL_X2 FILLER_0_43_285 ();
 FILLCELL_X1 FILLER_0_43_292 ();
 FILLCELL_X4 FILLER_0_43_296 ();
 FILLCELL_X1 FILLER_0_43_303 ();
 FILLCELL_X1 FILLER_0_43_307 ();
 FILLCELL_X8 FILLER_0_43_323 ();
 FILLCELL_X2 FILLER_0_43_331 ();
 FILLCELL_X1 FILLER_0_43_333 ();
 FILLCELL_X1 FILLER_0_43_345 ();
 FILLCELL_X1 FILLER_0_43_350 ();
 FILLCELL_X4 FILLER_0_43_354 ();
 FILLCELL_X2 FILLER_0_43_358 ();
 FILLCELL_X2 FILLER_0_43_394 ();
 FILLCELL_X2 FILLER_0_43_405 ();
 FILLCELL_X1 FILLER_0_43_407 ();
 FILLCELL_X32 FILLER_0_44_1 ();
 FILLCELL_X32 FILLER_0_44_33 ();
 FILLCELL_X32 FILLER_0_44_65 ();
 FILLCELL_X32 FILLER_0_44_97 ();
 FILLCELL_X32 FILLER_0_44_129 ();
 FILLCELL_X32 FILLER_0_44_161 ();
 FILLCELL_X32 FILLER_0_44_193 ();
 FILLCELL_X16 FILLER_0_44_225 ();
 FILLCELL_X4 FILLER_0_44_253 ();
 FILLCELL_X1 FILLER_0_44_257 ();
 FILLCELL_X4 FILLER_0_44_265 ();
 FILLCELL_X2 FILLER_0_44_269 ();
 FILLCELL_X2 FILLER_0_44_274 ();
 FILLCELL_X1 FILLER_0_44_276 ();
 FILLCELL_X2 FILLER_0_44_287 ();
 FILLCELL_X1 FILLER_0_44_289 ();
 FILLCELL_X2 FILLER_0_44_294 ();
 FILLCELL_X2 FILLER_0_44_313 ();
 FILLCELL_X1 FILLER_0_44_315 ();
 FILLCELL_X2 FILLER_0_44_319 ();
 FILLCELL_X2 FILLER_0_44_327 ();
 FILLCELL_X4 FILLER_0_44_333 ();
 FILLCELL_X1 FILLER_0_44_337 ();
 FILLCELL_X4 FILLER_0_44_341 ();
 FILLCELL_X2 FILLER_0_44_348 ();
 FILLCELL_X1 FILLER_0_44_350 ();
 FILLCELL_X2 FILLER_0_44_354 ();
 FILLCELL_X1 FILLER_0_44_356 ();
 FILLCELL_X4 FILLER_0_44_360 ();
 FILLCELL_X1 FILLER_0_44_364 ();
 FILLCELL_X2 FILLER_0_44_367 ();
 FILLCELL_X1 FILLER_0_44_369 ();
 FILLCELL_X1 FILLER_0_44_378 ();
 FILLCELL_X8 FILLER_0_44_381 ();
 FILLCELL_X4 FILLER_0_44_389 ();
 FILLCELL_X1 FILLER_0_44_407 ();
 FILLCELL_X32 FILLER_0_45_1 ();
 FILLCELL_X32 FILLER_0_45_33 ();
 FILLCELL_X32 FILLER_0_45_65 ();
 FILLCELL_X32 FILLER_0_45_97 ();
 FILLCELL_X32 FILLER_0_45_129 ();
 FILLCELL_X32 FILLER_0_45_161 ();
 FILLCELL_X32 FILLER_0_45_193 ();
 FILLCELL_X16 FILLER_0_45_225 ();
 FILLCELL_X8 FILLER_0_45_241 ();
 FILLCELL_X2 FILLER_0_45_249 ();
 FILLCELL_X2 FILLER_0_45_260 ();
 FILLCELL_X1 FILLER_0_45_262 ();
 FILLCELL_X2 FILLER_0_45_286 ();
 FILLCELL_X2 FILLER_0_45_291 ();
 FILLCELL_X2 FILLER_0_45_297 ();
 FILLCELL_X1 FILLER_0_45_299 ();
 FILLCELL_X1 FILLER_0_45_303 ();
 FILLCELL_X2 FILLER_0_45_307 ();
 FILLCELL_X4 FILLER_0_45_325 ();
 FILLCELL_X2 FILLER_0_45_329 ();
 FILLCELL_X1 FILLER_0_45_331 ();
 FILLCELL_X4 FILLER_0_45_335 ();
 FILLCELL_X2 FILLER_0_45_346 ();
 FILLCELL_X4 FILLER_0_45_356 ();
 FILLCELL_X1 FILLER_0_45_360 ();
 FILLCELL_X1 FILLER_0_45_364 ();
 FILLCELL_X8 FILLER_0_45_385 ();
 FILLCELL_X2 FILLER_0_45_393 ();
 FILLCELL_X1 FILLER_0_45_401 ();
 FILLCELL_X2 FILLER_0_45_405 ();
 FILLCELL_X1 FILLER_0_45_407 ();
 FILLCELL_X32 FILLER_0_46_1 ();
 FILLCELL_X32 FILLER_0_46_33 ();
 FILLCELL_X32 FILLER_0_46_65 ();
 FILLCELL_X32 FILLER_0_46_97 ();
 FILLCELL_X32 FILLER_0_46_129 ();
 FILLCELL_X32 FILLER_0_46_161 ();
 FILLCELL_X32 FILLER_0_46_193 ();
 FILLCELL_X32 FILLER_0_46_225 ();
 FILLCELL_X16 FILLER_0_46_257 ();
 FILLCELL_X2 FILLER_0_46_273 ();
 FILLCELL_X1 FILLER_0_46_275 ();
 FILLCELL_X2 FILLER_0_46_289 ();
 FILLCELL_X2 FILLER_0_46_298 ();
 FILLCELL_X1 FILLER_0_46_300 ();
 FILLCELL_X16 FILLER_0_46_307 ();
 FILLCELL_X4 FILLER_0_46_323 ();
 FILLCELL_X2 FILLER_0_46_327 ();
 FILLCELL_X1 FILLER_0_46_329 ();
 FILLCELL_X4 FILLER_0_46_334 ();
 FILLCELL_X1 FILLER_0_46_338 ();
 FILLCELL_X1 FILLER_0_46_342 ();
 FILLCELL_X8 FILLER_0_46_347 ();
 FILLCELL_X4 FILLER_0_46_355 ();
 FILLCELL_X2 FILLER_0_46_359 ();
 FILLCELL_X1 FILLER_0_46_361 ();
 FILLCELL_X2 FILLER_0_46_364 ();
 FILLCELL_X1 FILLER_0_46_371 ();
 FILLCELL_X2 FILLER_0_46_397 ();
 FILLCELL_X2 FILLER_0_46_406 ();
 FILLCELL_X32 FILLER_0_47_1 ();
 FILLCELL_X32 FILLER_0_47_33 ();
 FILLCELL_X32 FILLER_0_47_65 ();
 FILLCELL_X32 FILLER_0_47_97 ();
 FILLCELL_X32 FILLER_0_47_129 ();
 FILLCELL_X32 FILLER_0_47_161 ();
 FILLCELL_X32 FILLER_0_47_193 ();
 FILLCELL_X32 FILLER_0_47_225 ();
 FILLCELL_X32 FILLER_0_47_257 ();
 FILLCELL_X32 FILLER_0_47_289 ();
 FILLCELL_X8 FILLER_0_47_321 ();
 FILLCELL_X4 FILLER_0_47_329 ();
 FILLCELL_X1 FILLER_0_47_343 ();
 FILLCELL_X2 FILLER_0_47_360 ();
 FILLCELL_X2 FILLER_0_47_372 ();
 FILLCELL_X2 FILLER_0_47_390 ();
 FILLCELL_X32 FILLER_0_48_1 ();
 FILLCELL_X32 FILLER_0_48_33 ();
 FILLCELL_X32 FILLER_0_48_65 ();
 FILLCELL_X32 FILLER_0_48_97 ();
 FILLCELL_X32 FILLER_0_48_129 ();
 FILLCELL_X32 FILLER_0_48_161 ();
 FILLCELL_X32 FILLER_0_48_193 ();
 FILLCELL_X32 FILLER_0_48_225 ();
 FILLCELL_X32 FILLER_0_48_257 ();
 FILLCELL_X32 FILLER_0_48_289 ();
 FILLCELL_X16 FILLER_0_48_321 ();
 FILLCELL_X2 FILLER_0_48_337 ();
 FILLCELL_X1 FILLER_0_48_339 ();
 FILLCELL_X8 FILLER_0_48_356 ();
 FILLCELL_X4 FILLER_0_48_364 ();
 FILLCELL_X2 FILLER_0_48_368 ();
 FILLCELL_X1 FILLER_0_48_370 ();
 FILLCELL_X2 FILLER_0_48_386 ();
 FILLCELL_X1 FILLER_0_48_404 ();
 FILLCELL_X32 FILLER_0_49_1 ();
 FILLCELL_X32 FILLER_0_49_33 ();
 FILLCELL_X32 FILLER_0_49_65 ();
 FILLCELL_X32 FILLER_0_49_97 ();
 FILLCELL_X32 FILLER_0_49_129 ();
 FILLCELL_X32 FILLER_0_49_161 ();
 FILLCELL_X32 FILLER_0_49_193 ();
 FILLCELL_X32 FILLER_0_49_225 ();
 FILLCELL_X32 FILLER_0_49_257 ();
 FILLCELL_X32 FILLER_0_49_289 ();
 FILLCELL_X8 FILLER_0_49_321 ();
 FILLCELL_X4 FILLER_0_49_329 ();
 FILLCELL_X2 FILLER_0_49_333 ();
 FILLCELL_X1 FILLER_0_49_335 ();
 FILLCELL_X2 FILLER_0_49_360 ();
 FILLCELL_X4 FILLER_0_49_369 ();
 FILLCELL_X2 FILLER_0_49_373 ();
 FILLCELL_X1 FILLER_0_49_404 ();
 FILLCELL_X32 FILLER_0_50_1 ();
 FILLCELL_X32 FILLER_0_50_33 ();
 FILLCELL_X32 FILLER_0_50_65 ();
 FILLCELL_X32 FILLER_0_50_97 ();
 FILLCELL_X32 FILLER_0_50_129 ();
 FILLCELL_X32 FILLER_0_50_161 ();
 FILLCELL_X32 FILLER_0_50_193 ();
 FILLCELL_X32 FILLER_0_50_225 ();
 FILLCELL_X32 FILLER_0_50_257 ();
 FILLCELL_X32 FILLER_0_50_289 ();
 FILLCELL_X16 FILLER_0_50_321 ();
 FILLCELL_X4 FILLER_0_50_337 ();
 FILLCELL_X2 FILLER_0_50_341 ();
 FILLCELL_X1 FILLER_0_50_349 ();
 FILLCELL_X8 FILLER_0_50_353 ();
 FILLCELL_X2 FILLER_0_50_361 ();
 FILLCELL_X16 FILLER_0_50_366 ();
 FILLCELL_X2 FILLER_0_50_382 ();
 FILLCELL_X1 FILLER_0_50_384 ();
 FILLCELL_X16 FILLER_0_50_388 ();
 FILLCELL_X4 FILLER_0_50_404 ();
 FILLCELL_X32 FILLER_0_51_1 ();
 FILLCELL_X32 FILLER_0_51_33 ();
 FILLCELL_X32 FILLER_0_51_65 ();
 FILLCELL_X32 FILLER_0_51_97 ();
 FILLCELL_X32 FILLER_0_51_129 ();
 FILLCELL_X32 FILLER_0_51_161 ();
 FILLCELL_X32 FILLER_0_51_193 ();
 FILLCELL_X32 FILLER_0_51_225 ();
 FILLCELL_X32 FILLER_0_51_257 ();
 FILLCELL_X32 FILLER_0_51_289 ();
 FILLCELL_X32 FILLER_0_51_321 ();
 FILLCELL_X32 FILLER_0_51_353 ();
 FILLCELL_X16 FILLER_0_51_385 ();
 FILLCELL_X4 FILLER_0_51_401 ();
 FILLCELL_X2 FILLER_0_51_405 ();
 FILLCELL_X1 FILLER_0_51_407 ();
 FILLCELL_X32 FILLER_0_52_1 ();
 FILLCELL_X32 FILLER_0_52_33 ();
 FILLCELL_X32 FILLER_0_52_65 ();
 FILLCELL_X32 FILLER_0_52_97 ();
 FILLCELL_X32 FILLER_0_52_129 ();
 FILLCELL_X32 FILLER_0_52_161 ();
 FILLCELL_X32 FILLER_0_52_193 ();
 FILLCELL_X32 FILLER_0_52_225 ();
 FILLCELL_X32 FILLER_0_52_257 ();
 FILLCELL_X32 FILLER_0_52_289 ();
 FILLCELL_X32 FILLER_0_52_321 ();
 FILLCELL_X32 FILLER_0_52_353 ();
 FILLCELL_X16 FILLER_0_52_385 ();
 FILLCELL_X4 FILLER_0_52_401 ();
 FILLCELL_X2 FILLER_0_52_405 ();
 FILLCELL_X1 FILLER_0_52_407 ();
 FILLCELL_X32 FILLER_0_53_1 ();
 FILLCELL_X32 FILLER_0_53_33 ();
 FILLCELL_X32 FILLER_0_53_65 ();
 FILLCELL_X32 FILLER_0_53_97 ();
 FILLCELL_X32 FILLER_0_53_129 ();
 FILLCELL_X32 FILLER_0_53_161 ();
 FILLCELL_X32 FILLER_0_53_193 ();
 FILLCELL_X32 FILLER_0_53_225 ();
 FILLCELL_X32 FILLER_0_53_257 ();
 FILLCELL_X32 FILLER_0_53_289 ();
 FILLCELL_X32 FILLER_0_53_321 ();
 FILLCELL_X32 FILLER_0_53_353 ();
 FILLCELL_X16 FILLER_0_53_385 ();
 FILLCELL_X4 FILLER_0_53_401 ();
 FILLCELL_X2 FILLER_0_53_405 ();
 FILLCELL_X1 FILLER_0_53_407 ();
 FILLCELL_X32 FILLER_0_54_1 ();
 FILLCELL_X32 FILLER_0_54_33 ();
 FILLCELL_X32 FILLER_0_54_65 ();
 FILLCELL_X32 FILLER_0_54_97 ();
 FILLCELL_X32 FILLER_0_54_129 ();
 FILLCELL_X32 FILLER_0_54_161 ();
 FILLCELL_X32 FILLER_0_54_193 ();
 FILLCELL_X32 FILLER_0_54_225 ();
 FILLCELL_X32 FILLER_0_54_257 ();
 FILLCELL_X32 FILLER_0_54_289 ();
 FILLCELL_X16 FILLER_0_54_321 ();
 FILLCELL_X4 FILLER_0_54_337 ();
 FILLCELL_X2 FILLER_0_54_341 ();
 FILLCELL_X1 FILLER_0_54_343 ();
 FILLCELL_X2 FILLER_0_54_350 ();
 FILLCELL_X8 FILLER_0_54_355 ();
 FILLCELL_X4 FILLER_0_54_363 ();
 FILLCELL_X32 FILLER_0_54_370 ();
 FILLCELL_X4 FILLER_0_54_402 ();
 FILLCELL_X2 FILLER_0_54_406 ();
endmodule
