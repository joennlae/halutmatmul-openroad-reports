module fp_16_32_adder (operand_fp16_i,
    operand_fp32_i,
    result_o);
 input [15:0] operand_fp16_i;
 input [31:0] operand_fp32_i;
 output [31:0] result_o;

 wire net13;
 wire net3;
 wire net2;
 wire net1;
 wire \operand_fp16_fp32[13] ;
 wire \operand_fp16_fp32[14] ;
 wire \operand_fp16_fp32[15] ;
 wire \operand_fp16_fp32[16] ;
 wire \operand_fp16_fp32[17] ;
 wire \operand_fp16_fp32[18] ;
 wire \operand_fp16_fp32[19] ;
 wire net12;
 wire \operand_fp16_fp32[20] ;
 wire \operand_fp16_fp32[21] ;
 wire \operand_fp16_fp32[22] ;
 wire \operand_fp16_fp32[23] ;
 wire \operand_fp16_fp32[24] ;
 wire \operand_fp16_fp32[25] ;
 wire \operand_fp16_fp32[26] ;
 wire \operand_fp16_fp32[27] ;
 wire \operand_fp16_fp32[29] ;
 wire net11;
 wire net14;
 wire net10;
 wire net9;
 wire net8;
 wire net7;
 wire net6;
 wire net5;
 wire net4;
 wire \adder/_00_ ;
 wire \adder/_01_ ;
 wire \adder/_02_ ;
 wire \adder/_03_ ;
 wire \adder/_04_ ;
 wire \adder/_05_ ;
 wire \adder/_06_ ;
 wire \adder/_07_ ;
 wire \adder/_08_ ;
 wire \adder/_09_ ;
 wire \adder/_10_ ;
 wire \adder/_11_ ;
 wire \adder/_12_ ;
 wire \adder/_13_ ;
 wire \adder/_14_ ;
 wire \adder/_15_ ;
 wire \adder/_16_ ;
 wire \adder/_17_ ;
 wire \adder/_18_ ;
 wire \adder/_19_ ;
 wire \adder/exp_prenorm_d[0] ;
 wire \adder/exp_prenorm_d[1] ;
 wire \adder/exp_prenorm_d[2] ;
 wire \adder/exp_prenorm_d[3] ;
 wire \adder/exp_prenorm_d[4] ;
 wire \adder/exp_prenorm_d[5] ;
 wire \adder/exp_prenorm_d[6] ;
 wire \adder/exp_prenorm_d[7] ;
 wire net155;
 wire net154;
 wire \adder/hb_a_d ;
 wire \adder/hb_b_d ;
 wire \adder/mant_norm_d[23] ;
 wire net153;
 wire net143;
 wire net142;
 wire net141;
 wire net140;
 wire net139;
 wire net138;
 wire net137;
 wire net136;
 wire net135;
 wire net134;
 wire net152;
 wire \adder/mant_prenorm_d[20] ;
 wire \adder/mant_prenorm_d[21] ;
 wire \adder/mant_prenorm_d[22] ;
 wire \adder/mant_prenorm_d[23] ;
 wire \adder/mant_prenorm_d[24] ;
 wire \adder/mant_prenorm_d[25] ;
 wire \adder/mant_prenorm_d[26] ;
 wire \adder/mant_prenorm_d[27] ;
 wire \adder/mant_prenorm_d[28] ;
 wire \adder/mant_prenorm_d[29] ;
 wire net151;
 wire \adder/mant_prenorm_d[30] ;
 wire \adder/mant_prenorm_d[31] ;
 wire \adder/mant_prenorm_d[32] ;
 wire \adder/mant_prenorm_d[33] ;
 wire \adder/mant_prenorm_d[34] ;
 wire \adder/mant_prenorm_d[35] ;
 wire \adder/mant_prenorm_d[36] ;
 wire \adder/mant_prenorm_d[37] ;
 wire \adder/mant_prenorm_d[38] ;
 wire \adder/mant_prenorm_d[39] ;
 wire net150;
 wire \adder/mant_prenorm_d[40] ;
 wire \adder/mant_prenorm_d[41] ;
 wire \adder/mant_prenorm_d[42] ;
 wire \adder/mant_prenorm_d[43] ;
 wire \adder/mant_prenorm_d[44] ;
 wire \adder/mant_prenorm_d[45] ;
 wire \adder/mant_prenorm_d[46] ;
 wire \adder/mant_prenorm_d[47] ;
 wire net149;
 wire net148;
 wire net147;
 wire net146;
 wire net145;
 wire net144;
 wire net210;
 wire \adder/adder/_0000_ ;
 wire \adder/adder/_0001_ ;
 wire \adder/adder/_0002_ ;
 wire \adder/adder/_0003_ ;
 wire \adder/adder/_0004_ ;
 wire \adder/adder/_0005_ ;
 wire \adder/adder/_0006_ ;
 wire \adder/adder/_0007_ ;
 wire \adder/adder/_0008_ ;
 wire \adder/adder/_0009_ ;
 wire \adder/adder/_0010_ ;
 wire \adder/adder/_0011_ ;
 wire \adder/adder/_0012_ ;
 wire \adder/adder/_0013_ ;
 wire \adder/adder/_0014_ ;
 wire \adder/adder/_0015_ ;
 wire \adder/adder/_0016_ ;
 wire \adder/adder/_0017_ ;
 wire \adder/adder/_0018_ ;
 wire \adder/adder/_0019_ ;
 wire \adder/adder/_0020_ ;
 wire \adder/adder/_0021_ ;
 wire \adder/adder/_0022_ ;
 wire \adder/adder/_0023_ ;
 wire \adder/adder/_0024_ ;
 wire \adder/adder/_0025_ ;
 wire \adder/adder/_0026_ ;
 wire \adder/adder/_0027_ ;
 wire \adder/adder/_0028_ ;
 wire \adder/adder/_0029_ ;
 wire \adder/adder/_0030_ ;
 wire \adder/adder/_0031_ ;
 wire \adder/adder/_0032_ ;
 wire \adder/adder/_0033_ ;
 wire \adder/adder/_0034_ ;
 wire \adder/adder/_0035_ ;
 wire \adder/adder/_0036_ ;
 wire \adder/adder/_0037_ ;
 wire \adder/adder/_0038_ ;
 wire \adder/adder/_0039_ ;
 wire \adder/adder/_0040_ ;
 wire \adder/adder/_0041_ ;
 wire \adder/adder/_0042_ ;
 wire \adder/adder/_0043_ ;
 wire \adder/adder/_0044_ ;
 wire \adder/adder/_0045_ ;
 wire \adder/adder/_0046_ ;
 wire \adder/adder/_0047_ ;
 wire \adder/adder/_0048_ ;
 wire \adder/adder/_0049_ ;
 wire \adder/adder/_0050_ ;
 wire \adder/adder/_0051_ ;
 wire \adder/adder/_0052_ ;
 wire \adder/adder/_0053_ ;
 wire \adder/adder/_0054_ ;
 wire \adder/adder/_0055_ ;
 wire \adder/adder/_0056_ ;
 wire \adder/adder/_0057_ ;
 wire \adder/adder/_0058_ ;
 wire \adder/adder/_0059_ ;
 wire \adder/adder/_0060_ ;
 wire \adder/adder/_0061_ ;
 wire \adder/adder/_0062_ ;
 wire \adder/adder/_0063_ ;
 wire \adder/adder/_0064_ ;
 wire \adder/adder/_0065_ ;
 wire \adder/adder/_0066_ ;
 wire \adder/adder/_0067_ ;
 wire \adder/adder/_0068_ ;
 wire \adder/adder/_0069_ ;
 wire \adder/adder/_0070_ ;
 wire \adder/adder/_0071_ ;
 wire \adder/adder/_0072_ ;
 wire \adder/adder/_0073_ ;
 wire \adder/adder/_0074_ ;
 wire \adder/adder/_0075_ ;
 wire net160;
 wire \adder/adder/_0077_ ;
 wire \adder/adder/_0078_ ;
 wire \adder/adder/_0079_ ;
 wire \adder/adder/_0080_ ;
 wire net159;
 wire \adder/adder/_0082_ ;
 wire \adder/adder/_0083_ ;
 wire \adder/adder/_0084_ ;
 wire \adder/adder/_0085_ ;
 wire \adder/adder/_0086_ ;
 wire \adder/adder/_0087_ ;
 wire \adder/adder/_0088_ ;
 wire \adder/adder/_0089_ ;
 wire \adder/adder/_0090_ ;
 wire \adder/adder/_0091_ ;
 wire \adder/adder/_0092_ ;
 wire \adder/adder/_0093_ ;
 wire \adder/adder/_0094_ ;
 wire \adder/adder/_0095_ ;
 wire \adder/adder/_0096_ ;
 wire \adder/adder/_0097_ ;
 wire \adder/adder/_0098_ ;
 wire \adder/adder/_0099_ ;
 wire \adder/adder/_0100_ ;
 wire \adder/adder/_0101_ ;
 wire \adder/adder/_0102_ ;
 wire \adder/adder/_0103_ ;
 wire \adder/adder/_0104_ ;
 wire \adder/adder/_0105_ ;
 wire \adder/adder/_0106_ ;
 wire \adder/adder/_0107_ ;
 wire \adder/adder/_0108_ ;
 wire \adder/adder/_0109_ ;
 wire \adder/adder/_0110_ ;
 wire \adder/adder/_0111_ ;
 wire \adder/adder/_0112_ ;
 wire \adder/adder/_0113_ ;
 wire \adder/adder/_0114_ ;
 wire \adder/adder/_0115_ ;
 wire \adder/adder/_0116_ ;
 wire \adder/adder/_0117_ ;
 wire \adder/adder/_0118_ ;
 wire \adder/adder/_0119_ ;
 wire \adder/adder/_0120_ ;
 wire \adder/adder/_0121_ ;
 wire \adder/adder/_0122_ ;
 wire \adder/adder/_0123_ ;
 wire \adder/adder/_0124_ ;
 wire \adder/adder/_0125_ ;
 wire \adder/adder/_0126_ ;
 wire \adder/adder/_0127_ ;
 wire \adder/adder/_0128_ ;
 wire \adder/adder/_0129_ ;
 wire \adder/adder/_0130_ ;
 wire \adder/adder/_0131_ ;
 wire \adder/adder/_0132_ ;
 wire \adder/adder/_0133_ ;
 wire \adder/adder/_0134_ ;
 wire \adder/adder/_0135_ ;
 wire \adder/adder/_0136_ ;
 wire \adder/adder/_0137_ ;
 wire \adder/adder/_0138_ ;
 wire \adder/adder/_0139_ ;
 wire \adder/adder/_0140_ ;
 wire \adder/adder/_0141_ ;
 wire \adder/adder/_0142_ ;
 wire \adder/adder/_0143_ ;
 wire \adder/adder/_0144_ ;
 wire \adder/adder/_0145_ ;
 wire \adder/adder/_0146_ ;
 wire \adder/adder/_0147_ ;
 wire \adder/adder/_0148_ ;
 wire \adder/adder/_0149_ ;
 wire \adder/adder/_0150_ ;
 wire \adder/adder/_0151_ ;
 wire \adder/adder/_0152_ ;
 wire \adder/adder/_0153_ ;
 wire \adder/adder/_0154_ ;
 wire \adder/adder/_0155_ ;
 wire \adder/adder/_0156_ ;
 wire \adder/adder/_0157_ ;
 wire \adder/adder/_0158_ ;
 wire \adder/adder/_0159_ ;
 wire \adder/adder/_0160_ ;
 wire \adder/adder/_0161_ ;
 wire \adder/adder/_0162_ ;
 wire \adder/adder/_0163_ ;
 wire \adder/adder/_0164_ ;
 wire \adder/adder/_0165_ ;
 wire \adder/adder/_0166_ ;
 wire \adder/adder/_0167_ ;
 wire \adder/adder/_0168_ ;
 wire \adder/adder/_0169_ ;
 wire \adder/adder/_0170_ ;
 wire \adder/adder/_0171_ ;
 wire \adder/adder/_0172_ ;
 wire \adder/adder/_0173_ ;
 wire \adder/adder/_0174_ ;
 wire \adder/adder/_0175_ ;
 wire \adder/adder/_0176_ ;
 wire \adder/adder/_0177_ ;
 wire \adder/adder/_0178_ ;
 wire \adder/adder/_0179_ ;
 wire \adder/adder/_0180_ ;
 wire \adder/adder/_0181_ ;
 wire \adder/adder/_0182_ ;
 wire \adder/adder/_0183_ ;
 wire \adder/adder/_0184_ ;
 wire \adder/adder/_0185_ ;
 wire \adder/adder/_0186_ ;
 wire \adder/adder/_0187_ ;
 wire \adder/adder/_0188_ ;
 wire \adder/adder/_0189_ ;
 wire \adder/adder/_0190_ ;
 wire \adder/adder/_0191_ ;
 wire \adder/adder/_0192_ ;
 wire \adder/adder/_0193_ ;
 wire \adder/adder/_0194_ ;
 wire \adder/adder/_0195_ ;
 wire \adder/adder/_0196_ ;
 wire \adder/adder/_0197_ ;
 wire \adder/adder/_0198_ ;
 wire \adder/adder/_0199_ ;
 wire \adder/adder/_0200_ ;
 wire \adder/adder/_0201_ ;
 wire \adder/adder/_0202_ ;
 wire \adder/adder/_0203_ ;
 wire \adder/adder/_0204_ ;
 wire \adder/adder/_0205_ ;
 wire \adder/adder/_0206_ ;
 wire \adder/adder/_0207_ ;
 wire \adder/adder/_0208_ ;
 wire \adder/adder/_0209_ ;
 wire \adder/adder/_0210_ ;
 wire \adder/adder/_0211_ ;
 wire \adder/adder/_0212_ ;
 wire \adder/adder/_0213_ ;
 wire \adder/adder/_0214_ ;
 wire \adder/adder/_0215_ ;
 wire \adder/adder/_0216_ ;
 wire \adder/adder/_0217_ ;
 wire \adder/adder/_0218_ ;
 wire \adder/adder/_0219_ ;
 wire \adder/adder/_0220_ ;
 wire \adder/adder/_0221_ ;
 wire \adder/adder/_0222_ ;
 wire \adder/adder/_0223_ ;
 wire \adder/adder/_0224_ ;
 wire \adder/adder/_0225_ ;
 wire \adder/adder/_0226_ ;
 wire \adder/adder/_0227_ ;
 wire \adder/adder/_0228_ ;
 wire \adder/adder/_0229_ ;
 wire \adder/adder/_0230_ ;
 wire \adder/adder/_0231_ ;
 wire \adder/adder/_0232_ ;
 wire \adder/adder/_0233_ ;
 wire \adder/adder/_0234_ ;
 wire \adder/adder/_0235_ ;
 wire \adder/adder/_0236_ ;
 wire \adder/adder/_0237_ ;
 wire \adder/adder/_0238_ ;
 wire \adder/adder/_0239_ ;
 wire \adder/adder/_0240_ ;
 wire \adder/adder/_0241_ ;
 wire \adder/adder/_0242_ ;
 wire \adder/adder/_0243_ ;
 wire \adder/adder/_0244_ ;
 wire \adder/adder/_0245_ ;
 wire \adder/adder/_0246_ ;
 wire \adder/adder/_0247_ ;
 wire \adder/adder/_0248_ ;
 wire \adder/adder/_0249_ ;
 wire \adder/adder/_0250_ ;
 wire \adder/adder/_0251_ ;
 wire \adder/adder/_0252_ ;
 wire \adder/adder/_0253_ ;
 wire \adder/adder/_0254_ ;
 wire \adder/adder/_0255_ ;
 wire \adder/adder/_0256_ ;
 wire \adder/adder/_0257_ ;
 wire \adder/adder/_0258_ ;
 wire net158;
 wire \adder/adder/_0260_ ;
 wire \adder/adder/_0261_ ;
 wire net157;
 wire \adder/adder/_0263_ ;
 wire \adder/adder/_0264_ ;
 wire \adder/adder/_0265_ ;
 wire \adder/adder/_0266_ ;
 wire \adder/adder/_0267_ ;
 wire \adder/adder/_0268_ ;
 wire \adder/adder/_0269_ ;
 wire \adder/adder/_0270_ ;
 wire \adder/adder/_0271_ ;
 wire \adder/adder/_0272_ ;
 wire \adder/adder/_0273_ ;
 wire \adder/adder/_0274_ ;
 wire \adder/adder/_0275_ ;
 wire \adder/adder/_0276_ ;
 wire \adder/adder/_0277_ ;
 wire \adder/adder/_0278_ ;
 wire \adder/adder/_0279_ ;
 wire \adder/adder/_0280_ ;
 wire \adder/adder/_0281_ ;
 wire \adder/adder/_0282_ ;
 wire \adder/adder/_0283_ ;
 wire \adder/adder/_0284_ ;
 wire \adder/adder/_0285_ ;
 wire \adder/adder/_0286_ ;
 wire \adder/adder/_0287_ ;
 wire \adder/adder/_0288_ ;
 wire \adder/adder/_0289_ ;
 wire \adder/adder/_0290_ ;
 wire \adder/adder/_0291_ ;
 wire \adder/adder/_0292_ ;
 wire \adder/adder/_0293_ ;
 wire \adder/adder/_0294_ ;
 wire \adder/adder/_0295_ ;
 wire \adder/adder/_0296_ ;
 wire \adder/adder/_0297_ ;
 wire \adder/adder/_0298_ ;
 wire \adder/adder/_0299_ ;
 wire net156;
 wire \adder/adder/_0301_ ;
 wire \adder/adder/_0302_ ;
 wire \adder/adder/_0303_ ;
 wire \adder/adder/_0304_ ;
 wire \adder/adder/_0305_ ;
 wire \adder/adder/_0306_ ;
 wire \adder/adder/_0307_ ;
 wire \adder/adder/_0308_ ;
 wire \adder/adder/_0309_ ;
 wire \adder/adder/_0310_ ;
 wire \adder/adder/_0311_ ;
 wire \adder/adder/_0312_ ;
 wire \adder/adder/_0313_ ;
 wire \adder/adder/_0314_ ;
 wire \adder/adder/_0315_ ;
 wire \adder/adder/_0316_ ;
 wire \adder/adder/_0317_ ;
 wire \adder/adder/_0318_ ;
 wire \adder/adder/_0319_ ;
 wire net209;
 wire \adder/adder/_0321_ ;
 wire \adder/adder/_0322_ ;
 wire \adder/adder/_0323_ ;
 wire \adder/adder/_0324_ ;
 wire \adder/adder/_0325_ ;
 wire \adder/adder/_0326_ ;
 wire \adder/adder/_0327_ ;
 wire \adder/adder/_0328_ ;
 wire \adder/adder/_0329_ ;
 wire \adder/adder/_0330_ ;
 wire \adder/adder/_0331_ ;
 wire \adder/adder/_0332_ ;
 wire \adder/adder/_0333_ ;
 wire \adder/adder/_0334_ ;
 wire \adder/adder/_0335_ ;
 wire \adder/adder/_0336_ ;
 wire \adder/adder/_0337_ ;
 wire \adder/adder/_0338_ ;
 wire \adder/adder/_0339_ ;
 wire \adder/adder/_0340_ ;
 wire \adder/adder/_0341_ ;
 wire \adder/adder/_0342_ ;
 wire \adder/adder/_0343_ ;
 wire \adder/adder/_0344_ ;
 wire \adder/adder/_0345_ ;
 wire \adder/adder/_0346_ ;
 wire \adder/adder/_0347_ ;
 wire \adder/adder/_0348_ ;
 wire \adder/adder/_0349_ ;
 wire \adder/adder/_0350_ ;
 wire \adder/adder/_0351_ ;
 wire \adder/adder/_0352_ ;
 wire \adder/adder/_0353_ ;
 wire \adder/adder/_0354_ ;
 wire \adder/adder/_0355_ ;
 wire \adder/adder/_0356_ ;
 wire \adder/adder/_0357_ ;
 wire \adder/adder/_0358_ ;
 wire \adder/adder/_0359_ ;
 wire \adder/adder/_0360_ ;
 wire \adder/adder/_0361_ ;
 wire \adder/adder/_0362_ ;
 wire \adder/adder/_0363_ ;
 wire \adder/adder/_0364_ ;
 wire \adder/adder/_0365_ ;
 wire \adder/adder/_0366_ ;
 wire \adder/adder/_0367_ ;
 wire \adder/adder/_0368_ ;
 wire \adder/adder/_0369_ ;
 wire \adder/adder/_0370_ ;
 wire \adder/adder/_0371_ ;
 wire \adder/adder/_0372_ ;
 wire \adder/adder/_0373_ ;
 wire \adder/adder/_0374_ ;
 wire \adder/adder/_0375_ ;
 wire \adder/adder/_0376_ ;
 wire \adder/adder/_0377_ ;
 wire \adder/adder/_0378_ ;
 wire \adder/adder/_0379_ ;
 wire \adder/adder/_0380_ ;
 wire \adder/adder/_0381_ ;
 wire \adder/adder/_0382_ ;
 wire \adder/adder/_0383_ ;
 wire \adder/adder/_0384_ ;
 wire \adder/adder/_0385_ ;
 wire \adder/adder/_0386_ ;
 wire \adder/adder/_0387_ ;
 wire \adder/adder/_0388_ ;
 wire \adder/adder/_0389_ ;
 wire \adder/adder/_0390_ ;
 wire \adder/adder/_0391_ ;
 wire \adder/adder/_0392_ ;
 wire \adder/adder/_0393_ ;
 wire \adder/adder/_0394_ ;
 wire \adder/adder/_0395_ ;
 wire \adder/adder/_0396_ ;
 wire \adder/adder/_0397_ ;
 wire \adder/adder/_0398_ ;
 wire \adder/adder/_0399_ ;
 wire \adder/adder/_0400_ ;
 wire \adder/adder/_0401_ ;
 wire \adder/adder/_0402_ ;
 wire \adder/adder/_0403_ ;
 wire \adder/adder/_0404_ ;
 wire \adder/adder/_0405_ ;
 wire \adder/adder/_0406_ ;
 wire \adder/adder/_0407_ ;
 wire \adder/adder/_0408_ ;
 wire \adder/adder/_0409_ ;
 wire \adder/adder/_0410_ ;
 wire \adder/adder/_0411_ ;
 wire \adder/adder/_0412_ ;
 wire \adder/adder/_0413_ ;
 wire \adder/adder/_0414_ ;
 wire \adder/adder/_0415_ ;
 wire \adder/adder/_0416_ ;
 wire \adder/adder/_0417_ ;
 wire \adder/adder/_0418_ ;
 wire \adder/adder/_0419_ ;
 wire \adder/adder/_0420_ ;
 wire \adder/adder/_0421_ ;
 wire net208;
 wire \adder/adder/_0423_ ;
 wire \adder/adder/_0424_ ;
 wire \adder/adder/_0425_ ;
 wire \adder/adder/_0426_ ;
 wire \adder/adder/_0427_ ;
 wire \adder/adder/_0428_ ;
 wire \adder/adder/_0429_ ;
 wire \adder/adder/_0430_ ;
 wire \adder/adder/_0431_ ;
 wire \adder/adder/_0432_ ;
 wire \adder/adder/_0433_ ;
 wire \adder/adder/_0434_ ;
 wire \adder/adder/_0435_ ;
 wire \adder/adder/_0436_ ;
 wire \adder/adder/_0437_ ;
 wire \adder/adder/_0438_ ;
 wire \adder/adder/_0439_ ;
 wire \adder/adder/_0440_ ;
 wire \adder/adder/_0441_ ;
 wire \adder/adder/_0442_ ;
 wire \adder/adder/_0443_ ;
 wire \adder/adder/_0444_ ;
 wire \adder/adder/_0445_ ;
 wire \adder/adder/_0446_ ;
 wire \adder/adder/_0447_ ;
 wire \adder/adder/_0448_ ;
 wire \adder/adder/_0449_ ;
 wire \adder/adder/_0450_ ;
 wire \adder/adder/_0451_ ;
 wire \adder/adder/_0452_ ;
 wire \adder/adder/_0453_ ;
 wire \adder/adder/_0454_ ;
 wire \adder/adder/_0455_ ;
 wire \adder/adder/_0456_ ;
 wire \adder/adder/_0457_ ;
 wire \adder/adder/_0458_ ;
 wire \adder/adder/_0459_ ;
 wire \adder/adder/_0460_ ;
 wire \adder/adder/_0461_ ;
 wire \adder/adder/_0462_ ;
 wire \adder/adder/_0463_ ;
 wire \adder/adder/_0464_ ;
 wire \adder/adder/_0465_ ;
 wire \adder/adder/_0466_ ;
 wire \adder/adder/_0467_ ;
 wire \adder/adder/_0468_ ;
 wire \adder/adder/_0469_ ;
 wire \adder/adder/_0470_ ;
 wire \adder/adder/_0471_ ;
 wire \adder/adder/_0472_ ;
 wire \adder/adder/_0473_ ;
 wire \adder/adder/_0474_ ;
 wire net207;
 wire \adder/adder/_0476_ ;
 wire \adder/adder/_0477_ ;
 wire net206;
 wire net205;
 wire net204;
 wire net203;
 wire net201;
 wire net200;
 wire net199;
 wire \adder/adder/_0485_ ;
 wire net198;
 wire \adder/adder/_0487_ ;
 wire \adder/adder/_0488_ ;
 wire \adder/adder/_0489_ ;
 wire \adder/adder/_0490_ ;
 wire \adder/adder/_0491_ ;
 wire \adder/adder/_0492_ ;
 wire \adder/adder/_0493_ ;
 wire \adder/adder/_0494_ ;
 wire \adder/adder/_0495_ ;
 wire \adder/adder/_0496_ ;
 wire \adder/adder/_0497_ ;
 wire \adder/adder/_0498_ ;
 wire \adder/adder/_0499_ ;
 wire \adder/adder/_0500_ ;
 wire \adder/adder/_0501_ ;
 wire \adder/adder/_0502_ ;
 wire \adder/adder/_0503_ ;
 wire \adder/adder/_0504_ ;
 wire \adder/adder/_0505_ ;
 wire \adder/adder/_0506_ ;
 wire net197;
 wire \adder/adder/_0508_ ;
 wire net196;
 wire \adder/adder/_0510_ ;
 wire \adder/adder/_0511_ ;
 wire net195;
 wire \adder/adder/_0513_ ;
 wire net194;
 wire net193;
 wire \adder/adder/_0516_ ;
 wire \adder/adder/_0517_ ;
 wire net192;
 wire \adder/adder/_0519_ ;
 wire \adder/adder/_0520_ ;
 wire \adder/adder/_0521_ ;
 wire net191;
 wire net190;
 wire \adder/adder/_0524_ ;
 wire \adder/adder/_0525_ ;
 wire net189;
 wire \adder/adder/_0527_ ;
 wire net188;
 wire \adder/adder/_0529_ ;
 wire \adder/adder/_0530_ ;
 wire \adder/adder/_0531_ ;
 wire \adder/adder/_0532_ ;
 wire net187;
 wire net186;
 wire \adder/adder/_0535_ ;
 wire \adder/adder/_0536_ ;
 wire \adder/adder/_0537_ ;
 wire \adder/adder/_0538_ ;
 wire \adder/adder/_0539_ ;
 wire \adder/adder/_0540_ ;
 wire \adder/adder/_0541_ ;
 wire \adder/adder/_0542_ ;
 wire \adder/adder/_0543_ ;
 wire \adder/adder/_0544_ ;
 wire \adder/adder/_0545_ ;
 wire \adder/adder/_0546_ ;
 wire \adder/adder/_0547_ ;
 wire \adder/adder/_0548_ ;
 wire \adder/adder/_0549_ ;
 wire \adder/adder/_0550_ ;
 wire \adder/adder/_0551_ ;
 wire \adder/adder/_0552_ ;
 wire \adder/adder/_0553_ ;
 wire net185;
 wire \adder/adder/_0555_ ;
 wire \adder/adder/_0556_ ;
 wire \adder/adder/_0557_ ;
 wire \adder/adder/_0558_ ;
 wire \adder/adder/_0559_ ;
 wire \adder/adder/_0560_ ;
 wire net184;
 wire \adder/adder/_0562_ ;
 wire \adder/adder/_0563_ ;
 wire \adder/adder/_0564_ ;
 wire net183;
 wire \adder/adder/_0566_ ;
 wire net182;
 wire \adder/adder/_0568_ ;
 wire \adder/adder/_0569_ ;
 wire \adder/adder/_0570_ ;
 wire \adder/adder/_0571_ ;
 wire \adder/adder/_0572_ ;
 wire \adder/adder/_0573_ ;
 wire \adder/adder/_0574_ ;
 wire \adder/adder/_0575_ ;
 wire \adder/adder/_0576_ ;
 wire \adder/adder/_0577_ ;
 wire \adder/adder/_0578_ ;
 wire \adder/adder/_0579_ ;
 wire \adder/adder/_0580_ ;
 wire \adder/adder/_0581_ ;
 wire \adder/adder/_0582_ ;
 wire \adder/adder/_0583_ ;
 wire \adder/adder/_0584_ ;
 wire \adder/adder/_0585_ ;
 wire \adder/adder/_0586_ ;
 wire \adder/adder/_0587_ ;
 wire \adder/adder/_0588_ ;
 wire \adder/adder/_0589_ ;
 wire \adder/adder/_0590_ ;
 wire \adder/adder/_0591_ ;
 wire \adder/adder/_0592_ ;
 wire \adder/adder/_0593_ ;
 wire \adder/adder/_0594_ ;
 wire \adder/adder/_0595_ ;
 wire \adder/adder/_0596_ ;
 wire \adder/adder/_0597_ ;
 wire \adder/adder/_0598_ ;
 wire \adder/adder/_0599_ ;
 wire \adder/adder/_0600_ ;
 wire \adder/adder/_0601_ ;
 wire \adder/adder/_0602_ ;
 wire \adder/adder/_0603_ ;
 wire \adder/adder/_0604_ ;
 wire \adder/adder/_0605_ ;
 wire \adder/adder/_0606_ ;
 wire \adder/adder/_0607_ ;
 wire \adder/adder/_0608_ ;
 wire \adder/adder/_0609_ ;
 wire \adder/adder/_0610_ ;
 wire \adder/adder/_0611_ ;
 wire \adder/adder/_0612_ ;
 wire \adder/adder/_0613_ ;
 wire \adder/adder/_0614_ ;
 wire \adder/adder/_0615_ ;
 wire \adder/adder/_0616_ ;
 wire \adder/adder/_0617_ ;
 wire \adder/adder/_0618_ ;
 wire \adder/adder/_0619_ ;
 wire \adder/adder/_0620_ ;
 wire \adder/adder/_0621_ ;
 wire \adder/adder/_0622_ ;
 wire \adder/adder/_0623_ ;
 wire \adder/adder/_0624_ ;
 wire \adder/adder/_0625_ ;
 wire \adder/adder/_0626_ ;
 wire \adder/adder/_0627_ ;
 wire \adder/adder/_0628_ ;
 wire \adder/adder/_0629_ ;
 wire \adder/adder/_0630_ ;
 wire \adder/adder/_0631_ ;
 wire \adder/adder/_0632_ ;
 wire \adder/adder/_0633_ ;
 wire \adder/adder/_0634_ ;
 wire \adder/adder/_0635_ ;
 wire \adder/adder/_0636_ ;
 wire net181;
 wire \adder/adder/_0638_ ;
 wire \adder/adder/_0639_ ;
 wire \adder/adder/_0640_ ;
 wire \adder/adder/_0641_ ;
 wire \adder/adder/_0642_ ;
 wire \adder/adder/_0643_ ;
 wire \adder/adder/_0644_ ;
 wire \adder/adder/_0645_ ;
 wire \adder/adder/_0646_ ;
 wire \adder/adder/_0647_ ;
 wire \adder/adder/_0648_ ;
 wire \adder/adder/_0649_ ;
 wire \adder/adder/_0650_ ;
 wire \adder/adder/_0651_ ;
 wire \adder/adder/_0652_ ;
 wire \adder/adder/_0653_ ;
 wire \adder/adder/_0654_ ;
 wire \adder/adder/_0655_ ;
 wire \adder/adder/_0656_ ;
 wire \adder/adder/_0657_ ;
 wire \adder/adder/_0658_ ;
 wire \adder/adder/_0659_ ;
 wire \adder/adder/_0660_ ;
 wire \adder/adder/_0661_ ;
 wire \adder/adder/_0662_ ;
 wire \adder/adder/_0663_ ;
 wire \adder/adder/_0664_ ;
 wire \adder/adder/_0665_ ;
 wire \adder/adder/_0666_ ;
 wire \adder/adder/_0667_ ;
 wire \adder/adder/_0668_ ;
 wire \adder/adder/_0669_ ;
 wire \adder/adder/_0670_ ;
 wire \adder/adder/_0671_ ;
 wire \adder/adder/_0672_ ;
 wire \adder/adder/_0673_ ;
 wire \adder/adder/_0674_ ;
 wire \adder/adder/_0675_ ;
 wire \adder/adder/_0676_ ;
 wire \adder/adder/_0677_ ;
 wire \adder/adder/_0678_ ;
 wire \adder/adder/_0679_ ;
 wire \adder/adder/_0680_ ;
 wire \adder/adder/_0681_ ;
 wire \adder/adder/_0682_ ;
 wire \adder/adder/_0683_ ;
 wire \adder/adder/_0684_ ;
 wire \adder/adder/_0685_ ;
 wire \adder/adder/_0686_ ;
 wire \adder/adder/_0687_ ;
 wire \adder/adder/_0688_ ;
 wire \adder/adder/_0689_ ;
 wire \adder/adder/_0690_ ;
 wire \adder/adder/_0691_ ;
 wire \adder/adder/_0692_ ;
 wire \adder/adder/_0693_ ;
 wire \adder/adder/_0694_ ;
 wire \adder/adder/_0695_ ;
 wire \adder/adder/_0696_ ;
 wire \adder/adder/_0697_ ;
 wire \adder/adder/_0698_ ;
 wire \adder/adder/_0699_ ;
 wire \adder/adder/_0700_ ;
 wire \adder/adder/_0701_ ;
 wire \adder/adder/_0702_ ;
 wire \adder/adder/_0703_ ;
 wire \adder/adder/_0704_ ;
 wire \adder/adder/_0705_ ;
 wire \adder/adder/_0706_ ;
 wire \adder/adder/_0707_ ;
 wire \adder/adder/_0708_ ;
 wire \adder/adder/_0709_ ;
 wire \adder/adder/_0710_ ;
 wire \adder/adder/_0711_ ;
 wire \adder/adder/_0712_ ;
 wire \adder/adder/_0713_ ;
 wire \adder/adder/_0714_ ;
 wire \adder/adder/_0715_ ;
 wire \adder/adder/_0716_ ;
 wire \adder/adder/_0717_ ;
 wire \adder/adder/_0718_ ;
 wire \adder/adder/_0719_ ;
 wire \adder/adder/_0720_ ;
 wire \adder/adder/_0721_ ;
 wire \adder/adder/_0722_ ;
 wire \adder/adder/_0723_ ;
 wire \adder/adder/_0724_ ;
 wire \adder/adder/_0725_ ;
 wire \adder/adder/_0726_ ;
 wire \adder/adder/_0727_ ;
 wire \adder/adder/_0728_ ;
 wire \adder/adder/_0729_ ;
 wire \adder/adder/_0730_ ;
 wire \adder/adder/_0731_ ;
 wire \adder/adder/_0732_ ;
 wire \adder/adder/_0733_ ;
 wire \adder/adder/_0734_ ;
 wire \adder/adder/_0735_ ;
 wire \adder/adder/_0736_ ;
 wire \adder/adder/_0737_ ;
 wire \adder/adder/_0738_ ;
 wire \adder/adder/_0739_ ;
 wire \adder/adder/_0740_ ;
 wire net180;
 wire \adder/adder/_0742_ ;
 wire \adder/adder/_0743_ ;
 wire \adder/adder/_0744_ ;
 wire \adder/adder/_0745_ ;
 wire \adder/adder/_0746_ ;
 wire \adder/adder/_0747_ ;
 wire \adder/adder/_0748_ ;
 wire \adder/adder/_0749_ ;
 wire \adder/adder/_0750_ ;
 wire \adder/adder/_0751_ ;
 wire \adder/adder/_0752_ ;
 wire \adder/adder/_0753_ ;
 wire net179;
 wire net178;
 wire net177;
 wire net176;
 wire net175;
 wire \adder/adder/_0759_ ;
 wire \adder/adder/_0760_ ;
 wire \adder/adder/_0761_ ;
 wire net174;
 wire \adder/adder/_0763_ ;
 wire \adder/adder/_0764_ ;
 wire \adder/adder/_0765_ ;
 wire \adder/adder/_0766_ ;
 wire \adder/adder/_0767_ ;
 wire net173;
 wire \adder/adder/_0769_ ;
 wire \adder/adder/_0770_ ;
 wire \adder/adder/_0771_ ;
 wire \adder/adder/_0772_ ;
 wire \adder/adder/_0773_ ;
 wire \adder/adder/_0774_ ;
 wire \adder/adder/_0775_ ;
 wire \adder/adder/_0776_ ;
 wire \adder/adder/_0777_ ;
 wire \adder/adder/_0778_ ;
 wire \adder/adder/_0779_ ;
 wire \adder/adder/_0780_ ;
 wire \adder/adder/_0781_ ;
 wire \adder/adder/_0782_ ;
 wire net172;
 wire \adder/adder/_0784_ ;
 wire \adder/adder/_0785_ ;
 wire \adder/adder/_0786_ ;
 wire \adder/adder/_0787_ ;
 wire \adder/adder/_0788_ ;
 wire \adder/adder/_0789_ ;
 wire \adder/adder/_0790_ ;
 wire \adder/adder/_0791_ ;
 wire \adder/adder/_0792_ ;
 wire \adder/adder/_0793_ ;
 wire \adder/adder/_0794_ ;
 wire \adder/adder/_0795_ ;
 wire \adder/adder/_0796_ ;
 wire \adder/adder/_0797_ ;
 wire net171;
 wire \adder/adder/_0799_ ;
 wire net170;
 wire \adder/adder/_0801_ ;
 wire \adder/adder/_0802_ ;
 wire \adder/adder/_0803_ ;
 wire net169;
 wire \adder/adder/_0805_ ;
 wire \adder/adder/_0806_ ;
 wire \adder/adder/_0807_ ;
 wire \adder/adder/_0808_ ;
 wire \adder/adder/_0809_ ;
 wire \adder/adder/_0810_ ;
 wire \adder/adder/_0811_ ;
 wire net168;
 wire \adder/adder/_0813_ ;
 wire \adder/adder/_0814_ ;
 wire \adder/adder/_0815_ ;
 wire \adder/adder/_0816_ ;
 wire \adder/adder/_0817_ ;
 wire \adder/adder/_0818_ ;
 wire \adder/adder/_0819_ ;
 wire \adder/adder/_0820_ ;
 wire \adder/adder/_0821_ ;
 wire \adder/adder/_0822_ ;
 wire \adder/adder/_0823_ ;
 wire \adder/adder/_0824_ ;
 wire \adder/adder/_0825_ ;
 wire \adder/adder/_0826_ ;
 wire net167;
 wire \adder/adder/_0828_ ;
 wire \adder/adder/_0829_ ;
 wire \adder/adder/_0830_ ;
 wire \adder/adder/_0831_ ;
 wire \adder/adder/_0832_ ;
 wire \adder/adder/_0833_ ;
 wire \adder/adder/_0834_ ;
 wire \adder/adder/_0835_ ;
 wire \adder/adder/_0836_ ;
 wire \adder/adder/_0837_ ;
 wire \adder/adder/_0838_ ;
 wire \adder/adder/_0839_ ;
 wire \adder/adder/_0840_ ;
 wire \adder/adder/_0841_ ;
 wire \adder/adder/_0842_ ;
 wire \adder/adder/_0843_ ;
 wire net166;
 wire \adder/adder/_0845_ ;
 wire \adder/adder/_0846_ ;
 wire \adder/adder/_0847_ ;
 wire \adder/adder/_0848_ ;
 wire \adder/adder/_0849_ ;
 wire \adder/adder/_0850_ ;
 wire \adder/adder/_0851_ ;
 wire \adder/adder/_0852_ ;
 wire \adder/adder/_0853_ ;
 wire \adder/adder/_0854_ ;
 wire \adder/adder/_0855_ ;
 wire \adder/adder/_0856_ ;
 wire \adder/adder/_0857_ ;
 wire \adder/adder/_0858_ ;
 wire \adder/adder/_0859_ ;
 wire \adder/adder/_0860_ ;
 wire \adder/adder/_0861_ ;
 wire \adder/adder/_0862_ ;
 wire \adder/adder/_0863_ ;
 wire \adder/adder/_0864_ ;
 wire net165;
 wire net164;
 wire \adder/adder/_0867_ ;
 wire \adder/adder/_0868_ ;
 wire \adder/adder/_0869_ ;
 wire \adder/adder/_0870_ ;
 wire \adder/adder/_0871_ ;
 wire \adder/adder/_0872_ ;
 wire \adder/adder/_0873_ ;
 wire net163;
 wire \adder/adder/_0875_ ;
 wire \adder/adder/_0876_ ;
 wire \adder/adder/_0877_ ;
 wire \adder/adder/_0878_ ;
 wire \adder/adder/_0879_ ;
 wire \adder/adder/_0880_ ;
 wire \adder/adder/_0881_ ;
 wire \adder/adder/_0882_ ;
 wire \adder/adder/_0883_ ;
 wire \adder/adder/_0884_ ;
 wire \adder/adder/_0885_ ;
 wire \adder/adder/_0886_ ;
 wire \adder/adder/_0887_ ;
 wire \adder/adder/_0888_ ;
 wire \adder/adder/_0889_ ;
 wire \adder/adder/_0890_ ;
 wire \adder/adder/_0891_ ;
 wire \adder/adder/_0892_ ;
 wire \adder/adder/_0893_ ;
 wire \adder/adder/_0894_ ;
 wire \adder/adder/_0895_ ;
 wire \adder/adder/_0896_ ;
 wire \adder/adder/_0897_ ;
 wire \adder/adder/_0898_ ;
 wire \adder/adder/_0899_ ;
 wire \adder/adder/_0900_ ;
 wire \adder/adder/_0901_ ;
 wire \adder/adder/_0902_ ;
 wire \adder/adder/_0903_ ;
 wire \adder/adder/_0904_ ;
 wire \adder/adder/_0905_ ;
 wire \adder/adder/_0906_ ;
 wire \adder/adder/_0907_ ;
 wire \adder/adder/_0908_ ;
 wire \adder/adder/_0909_ ;
 wire \adder/adder/_0910_ ;
 wire \adder/adder/_0911_ ;
 wire \adder/adder/_0912_ ;
 wire \adder/adder/_0913_ ;
 wire \adder/adder/_0914_ ;
 wire \adder/adder/_0915_ ;
 wire \adder/adder/_0916_ ;
 wire \adder/adder/_0917_ ;
 wire \adder/adder/_0918_ ;
 wire \adder/adder/_0919_ ;
 wire \adder/adder/_0920_ ;
 wire \adder/adder/_0921_ ;
 wire \adder/adder/_0922_ ;
 wire \adder/adder/_0923_ ;
 wire \adder/adder/_0924_ ;
 wire \adder/adder/_0925_ ;
 wire \adder/adder/_0926_ ;
 wire \adder/adder/_0927_ ;
 wire \adder/adder/_0928_ ;
 wire \adder/adder/_0929_ ;
 wire \adder/adder/_0930_ ;
 wire \adder/adder/_0931_ ;
 wire \adder/adder/_0932_ ;
 wire \adder/adder/_0933_ ;
 wire \adder/adder/_0934_ ;
 wire \adder/adder/_0935_ ;
 wire \adder/adder/_0936_ ;
 wire \adder/adder/_0937_ ;
 wire \adder/adder/_0938_ ;
 wire \adder/adder/_0939_ ;
 wire \adder/adder/_0940_ ;
 wire \adder/adder/_0941_ ;
 wire \adder/adder/_0942_ ;
 wire \adder/adder/_0943_ ;
 wire \adder/adder/_0944_ ;
 wire \adder/adder/_0945_ ;
 wire \adder/adder/_0946_ ;
 wire \adder/adder/_0947_ ;
 wire \adder/adder/_0948_ ;
 wire \adder/adder/_0949_ ;
 wire \adder/adder/_0950_ ;
 wire \adder/adder/_0951_ ;
 wire \adder/adder/_0952_ ;
 wire \adder/adder/_0953_ ;
 wire \adder/adder/_0954_ ;
 wire net162;
 wire \adder/adder/_0956_ ;
 wire \adder/adder/_0957_ ;
 wire \adder/adder/_0958_ ;
 wire \adder/adder/_0959_ ;
 wire \adder/adder/_0960_ ;
 wire \adder/adder/_0961_ ;
 wire \adder/adder/_0962_ ;
 wire \adder/adder/_0963_ ;
 wire \adder/adder/_0964_ ;
 wire \adder/adder/_0965_ ;
 wire \adder/adder/_0966_ ;
 wire \adder/adder/_0967_ ;
 wire \adder/adder/_0968_ ;
 wire \adder/adder/_0969_ ;
 wire \adder/adder/_0970_ ;
 wire \adder/adder/_0971_ ;
 wire \adder/adder/_0972_ ;
 wire \adder/adder/_0973_ ;
 wire \adder/adder/_0974_ ;
 wire \adder/adder/_0975_ ;
 wire \adder/adder/_0976_ ;
 wire \adder/adder/_0977_ ;
 wire \adder/adder/_0978_ ;
 wire \adder/adder/_0979_ ;
 wire \adder/adder/_0980_ ;
 wire \adder/adder/_0981_ ;
 wire \adder/adder/_0982_ ;
 wire \adder/adder/_0983_ ;
 wire \adder/adder/_0984_ ;
 wire \adder/adder/_0985_ ;
 wire \adder/adder/_0986_ ;
 wire \adder/adder/_0987_ ;
 wire \adder/adder/_0988_ ;
 wire \adder/adder/_0989_ ;
 wire \adder/adder/_0990_ ;
 wire \adder/adder/_0991_ ;
 wire \adder/adder/_0992_ ;
 wire \adder/adder/_0993_ ;
 wire \adder/adder/_0994_ ;
 wire \adder/adder/_0995_ ;
 wire \adder/adder/_0996_ ;
 wire \adder/adder/_0997_ ;
 wire \adder/adder/_0998_ ;
 wire \adder/adder/_0999_ ;
 wire \adder/adder/_1000_ ;
 wire \adder/adder/_1001_ ;
 wire \adder/adder/_1002_ ;
 wire \adder/adder/_1003_ ;
 wire \adder/adder/_1004_ ;
 wire \adder/adder/_1005_ ;
 wire \adder/adder/_1006_ ;
 wire \adder/adder/_1007_ ;
 wire \adder/adder/_1008_ ;
 wire \adder/adder/_1009_ ;
 wire \adder/adder/_1010_ ;
 wire \adder/adder/_1011_ ;
 wire \adder/adder/_1012_ ;
 wire \adder/adder/_1013_ ;
 wire \adder/adder/_1014_ ;
 wire \adder/adder/_1015_ ;
 wire \adder/adder/_1016_ ;
 wire \adder/adder/_1017_ ;
 wire \adder/adder/_1018_ ;
 wire \adder/adder/_1019_ ;
 wire \adder/adder/_1020_ ;
 wire \adder/adder/_1021_ ;
 wire \adder/adder/_1022_ ;
 wire \adder/adder/_1023_ ;
 wire \adder/adder/_1024_ ;
 wire \adder/adder/_1025_ ;
 wire \adder/adder/_1026_ ;
 wire \adder/adder/_1027_ ;
 wire \adder/adder/_1028_ ;
 wire \adder/adder/_1029_ ;
 wire \adder/adder/_1030_ ;
 wire \adder/adder/_1031_ ;
 wire \adder/adder/_1032_ ;
 wire \adder/adder/_1033_ ;
 wire \adder/adder/_1034_ ;
 wire \adder/adder/_1035_ ;
 wire \adder/adder/_1036_ ;
 wire \adder/adder/_1037_ ;
 wire \adder/adder/_1038_ ;
 wire \adder/adder/_1039_ ;
 wire \adder/adder/_1040_ ;
 wire \adder/adder/_1041_ ;
 wire \adder/adder/_1042_ ;
 wire \adder/adder/_1043_ ;
 wire \adder/adder/_1044_ ;
 wire \adder/adder/_1045_ ;
 wire \adder/adder/_1046_ ;
 wire \adder/adder/_1047_ ;
 wire \adder/adder/_1048_ ;
 wire \adder/adder/_1049_ ;
 wire \adder/adder/_1050_ ;
 wire \adder/adder/_1051_ ;
 wire \adder/adder/_1052_ ;
 wire \adder/adder/_1053_ ;
 wire \adder/adder/_1054_ ;
 wire \adder/adder/_1055_ ;
 wire \adder/adder/_1056_ ;
 wire \adder/adder/_1057_ ;
 wire \adder/adder/_1058_ ;
 wire \adder/adder/_1059_ ;
 wire \adder/adder/_1060_ ;
 wire \adder/adder/_1061_ ;
 wire \adder/adder/_1062_ ;
 wire \adder/adder/_1063_ ;
 wire \adder/adder/_1064_ ;
 wire \adder/adder/_1065_ ;
 wire net161;
 wire \adder/adder/_1067_ ;
 wire \adder/adder/_1068_ ;
 wire \adder/adder/_1069_ ;
 wire \adder/adder/_1070_ ;
 wire \adder/adder/_1071_ ;
 wire \adder/adder/_1072_ ;
 wire \adder/adder/_1073_ ;
 wire \adder/adder/_1074_ ;
 wire \adder/adder/_1075_ ;
 wire \adder/adder/_1076_ ;
 wire \adder/adder/_1077_ ;
 wire \adder/adder/_1078_ ;
 wire \adder/adder/_1079_ ;
 wire \adder/adder/_1080_ ;
 wire \adder/adder/_1081_ ;
 wire \adder/adder/_1082_ ;
 wire \adder/adder/_1083_ ;
 wire \adder/adder/_1084_ ;
 wire \adder/adder/_1085_ ;
 wire \adder/adder/_1086_ ;
 wire \adder/adder/_1087_ ;
 wire \adder/adder/_1088_ ;
 wire \adder/adder/_1089_ ;
 wire \adder/adder/_1090_ ;
 wire \adder/adder/_1091_ ;
 wire \adder/adder/_1092_ ;
 wire \adder/adder/_1093_ ;
 wire \adder/adder/_1094_ ;
 wire \adder/adder/_1095_ ;
 wire \adder/adder/_1096_ ;
 wire \adder/adder/_1097_ ;
 wire \adder/adder/_1098_ ;
 wire \adder/adder/_1099_ ;
 wire \adder/adder/_1100_ ;
 wire \adder/adder/_1101_ ;
 wire \adder/adder/_1102_ ;
 wire \adder/adder/_1103_ ;
 wire \adder/adder/_1104_ ;
 wire \adder/adder/_1105_ ;
 wire \adder/adder/_1106_ ;
 wire net202;
 wire \adder/norm/Mant_leadingOne_D[0] ;
 wire \adder/norm/Mant_leadingOne_D[1] ;
 wire \adder/norm/Mant_leadingOne_D[2] ;
 wire \adder/norm/Mant_leadingOne_D[3] ;
 wire \adder/norm/Mant_leadingOne_D[4] ;
 wire \adder/norm/Mant_leadingOne_D[5] ;
 wire \adder/norm/Mant_zero_S ;
 wire \adder/norm/_0000_ ;
 wire \adder/norm/_0001_ ;
 wire \adder/norm/_0002_ ;
 wire \adder/norm/_0003_ ;
 wire \adder/norm/_0004_ ;
 wire \adder/norm/_0005_ ;
 wire \adder/norm/_0006_ ;
 wire \adder/norm/_0007_ ;
 wire \adder/norm/_0008_ ;
 wire \adder/norm/_0009_ ;
 wire \adder/norm/_0010_ ;
 wire \adder/norm/_0011_ ;
 wire \adder/norm/_0012_ ;
 wire \adder/norm/_0013_ ;
 wire \adder/norm/_0014_ ;
 wire \adder/norm/_0015_ ;
 wire \adder/norm/_0016_ ;
 wire \adder/norm/_0017_ ;
 wire \adder/norm/_0018_ ;
 wire \adder/norm/_0019_ ;
 wire \adder/norm/_0020_ ;
 wire \adder/norm/_0021_ ;
 wire \adder/norm/_0022_ ;
 wire \adder/norm/_0023_ ;
 wire \adder/norm/_0024_ ;
 wire \adder/norm/_0025_ ;
 wire \adder/norm/_0026_ ;
 wire \adder/norm/_0027_ ;
 wire \adder/norm/_0028_ ;
 wire \adder/norm/_0029_ ;
 wire \adder/norm/_0030_ ;
 wire \adder/norm/_0031_ ;
 wire net133;
 wire \adder/norm/_0033_ ;
 wire \adder/norm/_0034_ ;
 wire \adder/norm/_0035_ ;
 wire \adder/norm/_0036_ ;
 wire \adder/norm/_0037_ ;
 wire \adder/norm/_0038_ ;
 wire \adder/norm/_0039_ ;
 wire \adder/norm/_0040_ ;
 wire \adder/norm/_0041_ ;
 wire \adder/norm/_0042_ ;
 wire \adder/norm/_0043_ ;
 wire \adder/norm/_0044_ ;
 wire \adder/norm/_0045_ ;
 wire \adder/norm/_0046_ ;
 wire \adder/norm/_0047_ ;
 wire \adder/norm/_0048_ ;
 wire \adder/norm/_0049_ ;
 wire \adder/norm/_0050_ ;
 wire \adder/norm/_0051_ ;
 wire \adder/norm/_0052_ ;
 wire \adder/norm/_0053_ ;
 wire \adder/norm/_0054_ ;
 wire \adder/norm/_0055_ ;
 wire \adder/norm/_0056_ ;
 wire \adder/norm/_0057_ ;
 wire \adder/norm/_0058_ ;
 wire \adder/norm/_0059_ ;
 wire \adder/norm/_0060_ ;
 wire \adder/norm/_0061_ ;
 wire \adder/norm/_0062_ ;
 wire \adder/norm/_0063_ ;
 wire \adder/norm/_0064_ ;
 wire \adder/norm/_0065_ ;
 wire \adder/norm/_0066_ ;
 wire \adder/norm/_0067_ ;
 wire \adder/norm/_0068_ ;
 wire \adder/norm/_0069_ ;
 wire \adder/norm/_0070_ ;
 wire \adder/norm/_0071_ ;
 wire \adder/norm/_0072_ ;
 wire \adder/norm/_0073_ ;
 wire \adder/norm/_0074_ ;
 wire \adder/norm/_0075_ ;
 wire \adder/norm/_0076_ ;
 wire \adder/norm/_0077_ ;
 wire \adder/norm/_0078_ ;
 wire \adder/norm/_0079_ ;
 wire \adder/norm/_0080_ ;
 wire \adder/norm/_0081_ ;
 wire \adder/norm/_0082_ ;
 wire \adder/norm/_0083_ ;
 wire \adder/norm/_0084_ ;
 wire net51;
 wire \adder/norm/_0086_ ;
 wire \adder/norm/_0087_ ;
 wire \adder/norm/_0088_ ;
 wire \adder/norm/_0089_ ;
 wire \adder/norm/_0090_ ;
 wire net50;
 wire \adder/norm/_0092_ ;
 wire net49;
 wire \adder/norm/_0094_ ;
 wire net48;
 wire \adder/norm/_0096_ ;
 wire \adder/norm/_0097_ ;
 wire \adder/norm/_0098_ ;
 wire net47;
 wire \adder/norm/_0100_ ;
 wire \adder/norm/_0101_ ;
 wire net46;
 wire \adder/norm/_0103_ ;
 wire net45;
 wire \adder/norm/_0105_ ;
 wire \adder/norm/_0106_ ;
 wire net44;
 wire net43;
 wire \adder/norm/_0109_ ;
 wire \adder/norm/_0110_ ;
 wire \adder/norm/_0111_ ;
 wire \adder/norm/_0112_ ;
 wire \adder/norm/_0113_ ;
 wire \adder/norm/_0114_ ;
 wire \adder/norm/_0115_ ;
 wire \adder/norm/_0116_ ;
 wire \adder/norm/_0117_ ;
 wire net42;
 wire \adder/norm/_0119_ ;
 wire net41;
 wire \adder/norm/_0121_ ;
 wire net40;
 wire \adder/norm/_0123_ ;
 wire \adder/norm/_0124_ ;
 wire net39;
 wire \adder/norm/_0126_ ;
 wire \adder/norm/_0127_ ;
 wire \adder/norm/_0128_ ;
 wire net38;
 wire \adder/norm/_0130_ ;
 wire \adder/norm/_0131_ ;
 wire \adder/norm/_0132_ ;
 wire \adder/norm/_0133_ ;
 wire \adder/norm/_0134_ ;
 wire net37;
 wire \adder/norm/_0136_ ;
 wire \adder/norm/_0137_ ;
 wire \adder/norm/_0138_ ;
 wire \adder/norm/_0139_ ;
 wire net36;
 wire \adder/norm/_0141_ ;
 wire \adder/norm/_0142_ ;
 wire net35;
 wire \adder/norm/_0144_ ;
 wire \adder/norm/_0145_ ;
 wire \adder/norm/_0146_ ;
 wire net34;
 wire net33;
 wire \adder/norm/_0149_ ;
 wire net32;
 wire \adder/norm/_0151_ ;
 wire \adder/norm/_0152_ ;
 wire net31;
 wire \adder/norm/_0154_ ;
 wire net30;
 wire \adder/norm/_0156_ ;
 wire \adder/norm/_0157_ ;
 wire \adder/norm/_0158_ ;
 wire \adder/norm/_0159_ ;
 wire \adder/norm/_0160_ ;
 wire \adder/norm/_0161_ ;
 wire \adder/norm/_0162_ ;
 wire net29;
 wire \adder/norm/_0164_ ;
 wire \adder/norm/_0165_ ;
 wire \adder/norm/_0166_ ;
 wire \adder/norm/_0167_ ;
 wire \adder/norm/_0168_ ;
 wire \adder/norm/_0169_ ;
 wire \adder/norm/_0170_ ;
 wire \adder/norm/_0171_ ;
 wire \adder/norm/_0172_ ;
 wire \adder/norm/_0173_ ;
 wire \adder/norm/_0174_ ;
 wire \adder/norm/_0175_ ;
 wire \adder/norm/_0176_ ;
 wire \adder/norm/_0177_ ;
 wire \adder/norm/_0178_ ;
 wire \adder/norm/_0179_ ;
 wire \adder/norm/_0180_ ;
 wire \adder/norm/_0181_ ;
 wire \adder/norm/_0182_ ;
 wire \adder/norm/_0183_ ;
 wire \adder/norm/_0184_ ;
 wire \adder/norm/_0185_ ;
 wire \adder/norm/_0186_ ;
 wire \adder/norm/_0187_ ;
 wire \adder/norm/_0188_ ;
 wire \adder/norm/_0189_ ;
 wire \adder/norm/_0190_ ;
 wire net28;
 wire \adder/norm/_0192_ ;
 wire \adder/norm/_0193_ ;
 wire net27;
 wire \adder/norm/_0195_ ;
 wire net26;
 wire \adder/norm/_0197_ ;
 wire \adder/norm/_0198_ ;
 wire \adder/norm/_0199_ ;
 wire \adder/norm/_0200_ ;
 wire \adder/norm/_0201_ ;
 wire \adder/norm/_0202_ ;
 wire \adder/norm/_0203_ ;
 wire \adder/norm/_0204_ ;
 wire \adder/norm/_0205_ ;
 wire \adder/norm/_0206_ ;
 wire \adder/norm/_0207_ ;
 wire \adder/norm/_0208_ ;
 wire \adder/norm/_0209_ ;
 wire \adder/norm/_0210_ ;
 wire \adder/norm/_0211_ ;
 wire \adder/norm/_0212_ ;
 wire \adder/norm/_0213_ ;
 wire \adder/norm/_0214_ ;
 wire \adder/norm/_0215_ ;
 wire \adder/norm/_0216_ ;
 wire \adder/norm/_0217_ ;
 wire \adder/norm/_0218_ ;
 wire \adder/norm/_0219_ ;
 wire \adder/norm/_0220_ ;
 wire \adder/norm/_0221_ ;
 wire \adder/norm/_0222_ ;
 wire \adder/norm/_0223_ ;
 wire \adder/norm/_0224_ ;
 wire \adder/norm/_0225_ ;
 wire \adder/norm/_0226_ ;
 wire \adder/norm/_0227_ ;
 wire \adder/norm/_0228_ ;
 wire \adder/norm/_0229_ ;
 wire \adder/norm/_0230_ ;
 wire \adder/norm/_0231_ ;
 wire \adder/norm/_0232_ ;
 wire \adder/norm/_0233_ ;
 wire \adder/norm/_0234_ ;
 wire \adder/norm/_0235_ ;
 wire \adder/norm/_0236_ ;
 wire \adder/norm/_0237_ ;
 wire \adder/norm/_0238_ ;
 wire \adder/norm/_0239_ ;
 wire \adder/norm/_0240_ ;
 wire \adder/norm/_0241_ ;
 wire net25;
 wire \adder/norm/_0243_ ;
 wire net132;
 wire \adder/norm/_0245_ ;
 wire \adder/norm/_0246_ ;
 wire \adder/norm/_0247_ ;
 wire \adder/norm/_0248_ ;
 wire \adder/norm/_0249_ ;
 wire \adder/norm/_0250_ ;
 wire \adder/norm/_0251_ ;
 wire \adder/norm/_0252_ ;
 wire \adder/norm/_0253_ ;
 wire \adder/norm/_0254_ ;
 wire \adder/norm/_0255_ ;
 wire \adder/norm/_0256_ ;
 wire \adder/norm/_0257_ ;
 wire \adder/norm/_0258_ ;
 wire \adder/norm/_0259_ ;
 wire \adder/norm/_0260_ ;
 wire \adder/norm/_0261_ ;
 wire \adder/norm/_0262_ ;
 wire \adder/norm/_0263_ ;
 wire \adder/norm/_0264_ ;
 wire \adder/norm/_0265_ ;
 wire net131;
 wire \adder/norm/_0267_ ;
 wire \adder/norm/_0268_ ;
 wire \adder/norm/_0269_ ;
 wire \adder/norm/_0270_ ;
 wire \adder/norm/_0271_ ;
 wire \adder/norm/_0272_ ;
 wire \adder/norm/_0273_ ;
 wire \adder/norm/_0274_ ;
 wire \adder/norm/_0275_ ;
 wire \adder/norm/_0276_ ;
 wire \adder/norm/_0277_ ;
 wire \adder/norm/_0278_ ;
 wire \adder/norm/_0279_ ;
 wire \adder/norm/_0280_ ;
 wire \adder/norm/_0281_ ;
 wire \adder/norm/_0282_ ;
 wire \adder/norm/_0283_ ;
 wire \adder/norm/_0284_ ;
 wire \adder/norm/_0285_ ;
 wire \adder/norm/_0286_ ;
 wire \adder/norm/_0287_ ;
 wire \adder/norm/_0288_ ;
 wire \adder/norm/_0289_ ;
 wire \adder/norm/_0290_ ;
 wire \adder/norm/_0291_ ;
 wire \adder/norm/_0292_ ;
 wire \adder/norm/_0293_ ;
 wire \adder/norm/_0294_ ;
 wire \adder/norm/_0295_ ;
 wire \adder/norm/_0296_ ;
 wire \adder/norm/_0297_ ;
 wire \adder/norm/_0298_ ;
 wire \adder/norm/_0299_ ;
 wire \adder/norm/_0300_ ;
 wire \adder/norm/_0301_ ;
 wire \adder/norm/_0302_ ;
 wire \adder/norm/_0303_ ;
 wire \adder/norm/_0304_ ;
 wire \adder/norm/_0305_ ;
 wire \adder/norm/_0306_ ;
 wire \adder/norm/_0307_ ;
 wire \adder/norm/_0308_ ;
 wire \adder/norm/_0309_ ;
 wire \adder/norm/_0310_ ;
 wire \adder/norm/_0311_ ;
 wire \adder/norm/_0312_ ;
 wire \adder/norm/_0313_ ;
 wire \adder/norm/_0314_ ;
 wire \adder/norm/_0315_ ;
 wire \adder/norm/_0316_ ;
 wire \adder/norm/_0317_ ;
 wire \adder/norm/_0318_ ;
 wire \adder/norm/_0319_ ;
 wire \adder/norm/_0320_ ;
 wire \adder/norm/_0321_ ;
 wire \adder/norm/_0322_ ;
 wire \adder/norm/_0323_ ;
 wire \adder/norm/_0324_ ;
 wire \adder/norm/_0325_ ;
 wire \adder/norm/_0326_ ;
 wire \adder/norm/_0327_ ;
 wire \adder/norm/_0328_ ;
 wire \adder/norm/_0329_ ;
 wire \adder/norm/_0330_ ;
 wire \adder/norm/_0331_ ;
 wire \adder/norm/_0332_ ;
 wire \adder/norm/_0333_ ;
 wire \adder/norm/_0334_ ;
 wire \adder/norm/_0335_ ;
 wire \adder/norm/_0336_ ;
 wire \adder/norm/_0337_ ;
 wire \adder/norm/_0338_ ;
 wire \adder/norm/_0339_ ;
 wire \adder/norm/_0340_ ;
 wire \adder/norm/_0341_ ;
 wire \adder/norm/_0342_ ;
 wire \adder/norm/_0343_ ;
 wire \adder/norm/_0344_ ;
 wire \adder/norm/_0345_ ;
 wire \adder/norm/_0346_ ;
 wire \adder/norm/_0347_ ;
 wire \adder/norm/_0348_ ;
 wire net24;
 wire \adder/norm/_0350_ ;
 wire \adder/norm/_0351_ ;
 wire \adder/norm/_0352_ ;
 wire \adder/norm/_0353_ ;
 wire \adder/norm/_0354_ ;
 wire \adder/norm/_0355_ ;
 wire \adder/norm/_0356_ ;
 wire \adder/norm/_0357_ ;
 wire \adder/norm/_0358_ ;
 wire \adder/norm/_0359_ ;
 wire \adder/norm/_0360_ ;
 wire \adder/norm/_0361_ ;
 wire \adder/norm/_0362_ ;
 wire \adder/norm/_0363_ ;
 wire \adder/norm/_0364_ ;
 wire \adder/norm/_0365_ ;
 wire \adder/norm/_0366_ ;
 wire \adder/norm/_0367_ ;
 wire \adder/norm/_0368_ ;
 wire \adder/norm/_0369_ ;
 wire \adder/norm/_0370_ ;
 wire \adder/norm/_0371_ ;
 wire \adder/norm/_0372_ ;
 wire \adder/norm/_0373_ ;
 wire \adder/norm/_0374_ ;
 wire \adder/norm/_0375_ ;
 wire \adder/norm/_0376_ ;
 wire \adder/norm/_0377_ ;
 wire \adder/norm/_0378_ ;
 wire \adder/norm/_0379_ ;
 wire \adder/norm/_0380_ ;
 wire \adder/norm/_0381_ ;
 wire \adder/norm/_0382_ ;
 wire \adder/norm/_0383_ ;
 wire \adder/norm/_0384_ ;
 wire \adder/norm/_0385_ ;
 wire \adder/norm/_0386_ ;
 wire \adder/norm/_0387_ ;
 wire \adder/norm/_0388_ ;
 wire \adder/norm/_0389_ ;
 wire \adder/norm/_0390_ ;
 wire \adder/norm/_0391_ ;
 wire \adder/norm/_0392_ ;
 wire \adder/norm/_0393_ ;
 wire \adder/norm/_0394_ ;
 wire \adder/norm/_0395_ ;
 wire \adder/norm/_0396_ ;
 wire \adder/norm/_0397_ ;
 wire \adder/norm/_0398_ ;
 wire \adder/norm/_0399_ ;
 wire \adder/norm/_0400_ ;
 wire \adder/norm/_0401_ ;
 wire \adder/norm/_0402_ ;
 wire \adder/norm/_0403_ ;
 wire \adder/norm/_0404_ ;
 wire \adder/norm/_0405_ ;
 wire \adder/norm/_0406_ ;
 wire \adder/norm/_0407_ ;
 wire \adder/norm/_0408_ ;
 wire net130;
 wire \adder/norm/_0410_ ;
 wire \adder/norm/_0411_ ;
 wire \adder/norm/_0412_ ;
 wire \adder/norm/_0413_ ;
 wire \adder/norm/_0414_ ;
 wire \adder/norm/_0415_ ;
 wire \adder/norm/_0416_ ;
 wire \adder/norm/_0417_ ;
 wire \adder/norm/_0418_ ;
 wire \adder/norm/_0419_ ;
 wire \adder/norm/_0420_ ;
 wire \adder/norm/_0421_ ;
 wire \adder/norm/_0422_ ;
 wire \adder/norm/_0423_ ;
 wire \adder/norm/_0424_ ;
 wire \adder/norm/_0425_ ;
 wire \adder/norm/_0426_ ;
 wire \adder/norm/_0427_ ;
 wire \adder/norm/_0428_ ;
 wire \adder/norm/_0429_ ;
 wire \adder/norm/_0430_ ;
 wire \adder/norm/_0431_ ;
 wire \adder/norm/_0432_ ;
 wire \adder/norm/_0433_ ;
 wire \adder/norm/_0434_ ;
 wire \adder/norm/_0435_ ;
 wire \adder/norm/_0436_ ;
 wire \adder/norm/_0437_ ;
 wire \adder/norm/_0438_ ;
 wire \adder/norm/_0439_ ;
 wire \adder/norm/_0440_ ;
 wire \adder/norm/_0441_ ;
 wire \adder/norm/_0442_ ;
 wire \adder/norm/_0443_ ;
 wire \adder/norm/_0444_ ;
 wire \adder/norm/_0445_ ;
 wire \adder/norm/_0446_ ;
 wire \adder/norm/_0447_ ;
 wire \adder/norm/_0448_ ;
 wire \adder/norm/_0449_ ;
 wire \adder/norm/_0450_ ;
 wire \adder/norm/_0451_ ;
 wire \adder/norm/_0452_ ;
 wire \adder/norm/_0453_ ;
 wire \adder/norm/_0454_ ;
 wire \adder/norm/_0455_ ;
 wire \adder/norm/_0456_ ;
 wire \adder/norm/_0457_ ;
 wire \adder/norm/_0458_ ;
 wire \adder/norm/_0459_ ;
 wire \adder/norm/_0460_ ;
 wire \adder/norm/_0461_ ;
 wire \adder/norm/_0462_ ;
 wire \adder/norm/_0463_ ;
 wire \adder/norm/_0464_ ;
 wire \adder/norm/_0465_ ;
 wire \adder/norm/_0466_ ;
 wire \adder/norm/_0467_ ;
 wire \adder/norm/_0468_ ;
 wire \adder/norm/_0469_ ;
 wire \adder/norm/_0470_ ;
 wire \adder/norm/_0471_ ;
 wire \adder/norm/_0472_ ;
 wire \adder/norm/_0473_ ;
 wire \adder/norm/_0474_ ;
 wire \adder/norm/_0475_ ;
 wire \adder/norm/_0476_ ;
 wire \adder/norm/_0477_ ;
 wire \adder/norm/_0478_ ;
 wire \adder/norm/_0479_ ;
 wire \adder/norm/_0480_ ;
 wire \adder/norm/_0481_ ;
 wire \adder/norm/_0482_ ;
 wire \adder/norm/_0483_ ;
 wire \adder/norm/_0484_ ;
 wire \adder/norm/_0485_ ;
 wire \adder/norm/_0486_ ;
 wire \adder/norm/_0487_ ;
 wire \adder/norm/_0488_ ;
 wire \adder/norm/_0489_ ;
 wire \adder/norm/_0490_ ;
 wire \adder/norm/_0491_ ;
 wire \adder/norm/_0492_ ;
 wire \adder/norm/_0493_ ;
 wire \adder/norm/_0494_ ;
 wire \adder/norm/_0495_ ;
 wire \adder/norm/_0496_ ;
 wire \adder/norm/_0497_ ;
 wire \adder/norm/_0498_ ;
 wire \adder/norm/_0499_ ;
 wire \adder/norm/_0500_ ;
 wire \adder/norm/_0501_ ;
 wire \adder/norm/_0502_ ;
 wire \adder/norm/_0503_ ;
 wire \adder/norm/_0504_ ;
 wire \adder/norm/_0505_ ;
 wire \adder/norm/_0506_ ;
 wire \adder/norm/_0507_ ;
 wire \adder/norm/_0508_ ;
 wire \adder/norm/_0509_ ;
 wire \adder/norm/_0510_ ;
 wire \adder/norm/_0511_ ;
 wire \adder/norm/_0512_ ;
 wire \adder/norm/_0513_ ;
 wire \adder/norm/_0514_ ;
 wire \adder/norm/_0515_ ;
 wire \adder/norm/_0516_ ;
 wire \adder/norm/_0517_ ;
 wire \adder/norm/_0518_ ;
 wire \adder/norm/_0519_ ;
 wire \adder/norm/_0520_ ;
 wire \adder/norm/_0521_ ;
 wire \adder/norm/_0522_ ;
 wire \adder/norm/_0523_ ;
 wire \adder/norm/_0524_ ;
 wire \adder/norm/_0525_ ;
 wire \adder/norm/_0526_ ;
 wire \adder/norm/_0527_ ;
 wire \adder/norm/_0528_ ;
 wire \adder/norm/_0529_ ;
 wire \adder/norm/_0530_ ;
 wire \adder/norm/_0531_ ;
 wire \adder/norm/_0532_ ;
 wire \adder/norm/_0533_ ;
 wire \adder/norm/_0534_ ;
 wire \adder/norm/_0535_ ;
 wire \adder/norm/_0536_ ;
 wire \adder/norm/_0537_ ;
 wire \adder/norm/_0538_ ;
 wire \adder/norm/_0539_ ;
 wire \adder/norm/_0540_ ;
 wire \adder/norm/_0541_ ;
 wire \adder/norm/_0542_ ;
 wire \adder/norm/_0543_ ;
 wire \adder/norm/_0544_ ;
 wire \adder/norm/_0545_ ;
 wire \adder/norm/_0546_ ;
 wire \adder/norm/_0547_ ;
 wire \adder/norm/_0548_ ;
 wire \adder/norm/_0549_ ;
 wire \adder/norm/_0550_ ;
 wire \adder/norm/_0551_ ;
 wire \adder/norm/_0552_ ;
 wire \adder/norm/_0553_ ;
 wire \adder/norm/_0554_ ;
 wire \adder/norm/_0555_ ;
 wire \adder/norm/_0556_ ;
 wire \adder/norm/_0557_ ;
 wire \adder/norm/_0558_ ;
 wire \adder/norm/_0559_ ;
 wire \adder/norm/_0560_ ;
 wire \adder/norm/_0561_ ;
 wire \adder/norm/_0562_ ;
 wire \adder/norm/_0563_ ;
 wire \adder/norm/_0564_ ;
 wire \adder/norm/_0565_ ;
 wire \adder/norm/_0566_ ;
 wire \adder/norm/_0567_ ;
 wire \adder/norm/_0568_ ;
 wire \adder/norm/_0569_ ;
 wire \adder/norm/_0570_ ;
 wire \adder/norm/_0571_ ;
 wire \adder/norm/_0572_ ;
 wire \adder/norm/_0573_ ;
 wire \adder/norm/_0574_ ;
 wire \adder/norm/_0575_ ;
 wire \adder/norm/_0576_ ;
 wire \adder/norm/_0577_ ;
 wire \adder/norm/_0578_ ;
 wire \adder/norm/_0579_ ;
 wire \adder/norm/_0580_ ;
 wire \adder/norm/_0581_ ;
 wire \adder/norm/_0582_ ;
 wire \adder/norm/_0583_ ;
 wire \adder/norm/_0584_ ;
 wire \adder/norm/_0585_ ;
 wire \adder/norm/_0586_ ;
 wire \adder/norm/_0587_ ;
 wire \adder/norm/_0588_ ;
 wire \adder/norm/_0589_ ;
 wire \adder/norm/_0590_ ;
 wire \adder/norm/_0591_ ;
 wire \adder/norm/_0592_ ;
 wire \adder/norm/_0593_ ;
 wire \adder/norm/_0594_ ;
 wire \adder/norm/_0595_ ;
 wire \adder/norm/_0596_ ;
 wire \adder/norm/_0597_ ;
 wire \adder/norm/_0598_ ;
 wire \adder/norm/_0599_ ;
 wire \adder/norm/_0600_ ;
 wire \adder/norm/_0601_ ;
 wire \adder/norm/_0602_ ;
 wire \adder/norm/_0603_ ;
 wire \adder/norm/_0604_ ;
 wire \adder/norm/_0605_ ;
 wire \adder/norm/_0606_ ;
 wire \adder/norm/_0607_ ;
 wire \adder/norm/_0608_ ;
 wire \adder/norm/_0609_ ;
 wire \adder/norm/_0610_ ;
 wire \adder/norm/_0611_ ;
 wire \adder/norm/_0612_ ;
 wire \adder/norm/_0613_ ;
 wire \adder/norm/_0614_ ;
 wire \adder/norm/_0615_ ;
 wire \adder/norm/_0616_ ;
 wire \adder/norm/_0617_ ;
 wire \adder/norm/_0618_ ;
 wire \adder/norm/_0619_ ;
 wire \adder/norm/_0620_ ;
 wire \adder/norm/_0621_ ;
 wire \adder/norm/_0622_ ;
 wire \adder/norm/_0623_ ;
 wire \adder/norm/_0624_ ;
 wire \adder/norm/_0625_ ;
 wire \adder/norm/_0626_ ;
 wire \adder/norm/_0627_ ;
 wire \adder/norm/_0628_ ;
 wire \adder/norm/_0629_ ;
 wire \adder/norm/_0630_ ;
 wire \adder/norm/_0631_ ;
 wire \adder/norm/_0632_ ;
 wire \adder/norm/_0633_ ;
 wire \adder/norm/_0634_ ;
 wire \adder/norm/_0635_ ;
 wire \adder/norm/_0636_ ;
 wire \adder/norm/_0637_ ;
 wire \adder/norm/_0638_ ;
 wire net129;
 wire \adder/norm/_0640_ ;
 wire \adder/norm/_0641_ ;
 wire \adder/norm/_0642_ ;
 wire \adder/norm/_0643_ ;
 wire \adder/norm/_0644_ ;
 wire \adder/norm/_0645_ ;
 wire \adder/norm/_0646_ ;
 wire \adder/norm/_0647_ ;
 wire \adder/norm/_0648_ ;
 wire \adder/norm/_0649_ ;
 wire \adder/norm/_0650_ ;
 wire \adder/norm/_0651_ ;
 wire \adder/norm/_0652_ ;
 wire \adder/norm/_0653_ ;
 wire \adder/norm/_0654_ ;
 wire \adder/norm/_0655_ ;
 wire \adder/norm/_0656_ ;
 wire \adder/norm/_0657_ ;
 wire \adder/norm/_0658_ ;
 wire \adder/norm/_0659_ ;
 wire \adder/norm/_0660_ ;
 wire net128;
 wire \adder/norm/_0662_ ;
 wire \adder/norm/_0663_ ;
 wire \adder/norm/_0664_ ;
 wire \adder/norm/_0665_ ;
 wire \adder/norm/_0666_ ;
 wire \adder/norm/_0667_ ;
 wire \adder/norm/_0668_ ;
 wire \adder/norm/_0669_ ;
 wire \adder/norm/_0670_ ;
 wire net127;
 wire \adder/norm/_0672_ ;
 wire \adder/norm/_0673_ ;
 wire net126;
 wire net125;
 wire \adder/norm/_0676_ ;
 wire \adder/norm/_0677_ ;
 wire \adder/norm/_0678_ ;
 wire \adder/norm/_0679_ ;
 wire \adder/norm/_0680_ ;
 wire \adder/norm/_0681_ ;
 wire net124;
 wire net123;
 wire \adder/norm/_0684_ ;
 wire net122;
 wire net121;
 wire net120;
 wire \adder/norm/_0688_ ;
 wire net119;
 wire net118;
 wire \adder/norm/_0691_ ;
 wire net117;
 wire \adder/norm/_0693_ ;
 wire \adder/norm/_0694_ ;
 wire net116;
 wire \adder/norm/_0696_ ;
 wire net115;
 wire \adder/norm/_0698_ ;
 wire \adder/norm/_0699_ ;
 wire net114;
 wire \adder/norm/_0701_ ;
 wire \adder/norm/_0702_ ;
 wire \adder/norm/_0703_ ;
 wire net113;
 wire \adder/norm/_0705_ ;
 wire net112;
 wire net111;
 wire net110;
 wire \adder/norm/_0709_ ;
 wire \adder/norm/_0710_ ;
 wire net109;
 wire \adder/norm/_0712_ ;
 wire \adder/norm/_0713_ ;
 wire \adder/norm/_0714_ ;
 wire \adder/norm/_0715_ ;
 wire \adder/norm/_0716_ ;
 wire \adder/norm/_0717_ ;
 wire net108;
 wire net107;
 wire \adder/norm/_0720_ ;
 wire net106;
 wire \adder/norm/_0722_ ;
 wire \adder/norm/_0723_ ;
 wire net105;
 wire \adder/norm/_0725_ ;
 wire \adder/norm/_0726_ ;
 wire \adder/norm/_0727_ ;
 wire \adder/norm/_0728_ ;
 wire net104;
 wire \adder/norm/_0730_ ;
 wire \adder/norm/_0731_ ;
 wire \adder/norm/_0732_ ;
 wire \adder/norm/_0733_ ;
 wire net103;
 wire \adder/norm/_0735_ ;
 wire net102;
 wire \adder/norm/_0737_ ;
 wire \adder/norm/_0738_ ;
 wire \adder/norm/_0739_ ;
 wire \adder/norm/_0740_ ;
 wire \adder/norm/_0741_ ;
 wire \adder/norm/_0742_ ;
 wire \adder/norm/_0743_ ;
 wire net101;
 wire \adder/norm/_0745_ ;
 wire \adder/norm/_0746_ ;
 wire \adder/norm/_0747_ ;
 wire net100;
 wire net99;
 wire \adder/norm/_0750_ ;
 wire \adder/norm/_0751_ ;
 wire \adder/norm/_0752_ ;
 wire \adder/norm/_0753_ ;
 wire \adder/norm/_0754_ ;
 wire \adder/norm/_0755_ ;
 wire \adder/norm/_0756_ ;
 wire \adder/norm/_0757_ ;
 wire \adder/norm/_0758_ ;
 wire \adder/norm/_0759_ ;
 wire \adder/norm/_0760_ ;
 wire \adder/norm/_0761_ ;
 wire net98;
 wire net97;
 wire \adder/norm/_0764_ ;
 wire \adder/norm/_0765_ ;
 wire net96;
 wire net95;
 wire \adder/norm/_0768_ ;
 wire net94;
 wire \adder/norm/_0770_ ;
 wire \adder/norm/_0771_ ;
 wire \adder/norm/_0772_ ;
 wire net93;
 wire \adder/norm/_0774_ ;
 wire \adder/norm/_0775_ ;
 wire \adder/norm/_0776_ ;
 wire \adder/norm/_0777_ ;
 wire \adder/norm/_0778_ ;
 wire \adder/norm/_0779_ ;
 wire net92;
 wire net91;
 wire \adder/norm/_0782_ ;
 wire \adder/norm/_0783_ ;
 wire \adder/norm/_0784_ ;
 wire \adder/norm/_0785_ ;
 wire \adder/norm/_0786_ ;
 wire \adder/norm/_0787_ ;
 wire \adder/norm/_0788_ ;
 wire \adder/norm/_0789_ ;
 wire \adder/norm/_0790_ ;
 wire net90;
 wire \adder/norm/_0792_ ;
 wire \adder/norm/_0793_ ;
 wire net89;
 wire \adder/norm/_0795_ ;
 wire \adder/norm/_0796_ ;
 wire \adder/norm/_0797_ ;
 wire \adder/norm/_0798_ ;
 wire \adder/norm/_0799_ ;
 wire \adder/norm/_0800_ ;
 wire \adder/norm/_0801_ ;
 wire \adder/norm/_0802_ ;
 wire \adder/norm/_0803_ ;
 wire net88;
 wire net87;
 wire \adder/norm/_0806_ ;
 wire \adder/norm/_0807_ ;
 wire \adder/norm/_0808_ ;
 wire \adder/norm/_0809_ ;
 wire \adder/norm/_0810_ ;
 wire \adder/norm/_0811_ ;
 wire \adder/norm/_0812_ ;
 wire \adder/norm/_0813_ ;
 wire \adder/norm/_0814_ ;
 wire \adder/norm/_0815_ ;
 wire \adder/norm/_0816_ ;
 wire \adder/norm/_0817_ ;
 wire \adder/norm/_0818_ ;
 wire \adder/norm/_0819_ ;
 wire \adder/norm/_0820_ ;
 wire net86;
 wire net85;
 wire \adder/norm/_0823_ ;
 wire \adder/norm/_0824_ ;
 wire \adder/norm/_0825_ ;
 wire \adder/norm/_0826_ ;
 wire \adder/norm/_0827_ ;
 wire \adder/norm/_0828_ ;
 wire \adder/norm/_0829_ ;
 wire net84;
 wire net83;
 wire net82;
 wire net81;
 wire \adder/norm/_0834_ ;
 wire \adder/norm/_0835_ ;
 wire \adder/norm/_0836_ ;
 wire net80;
 wire \adder/norm/_0838_ ;
 wire \adder/norm/_0839_ ;
 wire \adder/norm/_0840_ ;
 wire \adder/norm/_0841_ ;
 wire net79;
 wire net78;
 wire net77;
 wire \adder/norm/_0845_ ;
 wire net76;
 wire \adder/norm/_0847_ ;
 wire \adder/norm/_0848_ ;
 wire net75;
 wire \adder/norm/_0850_ ;
 wire \adder/norm/_0851_ ;
 wire \adder/norm/_0852_ ;
 wire \adder/norm/_0853_ ;
 wire \adder/norm/_0854_ ;
 wire \adder/norm/_0855_ ;
 wire net74;
 wire \adder/norm/_0857_ ;
 wire \adder/norm/_0858_ ;
 wire net73;
 wire \adder/norm/_0860_ ;
 wire \adder/norm/_0861_ ;
 wire net72;
 wire \adder/norm/_0863_ ;
 wire \adder/norm/_0864_ ;
 wire net71;
 wire net70;
 wire \adder/norm/_0867_ ;
 wire \adder/norm/_0868_ ;
 wire \adder/norm/_0869_ ;
 wire \adder/norm/_0870_ ;
 wire net69;
 wire \adder/norm/_0872_ ;
 wire \adder/norm/_0873_ ;
 wire \adder/norm/_0874_ ;
 wire \adder/norm/_0875_ ;
 wire \adder/norm/_0876_ ;
 wire \adder/norm/_0877_ ;
 wire \adder/norm/_0878_ ;
 wire \adder/norm/_0879_ ;
 wire net68;
 wire \adder/norm/_0881_ ;
 wire \adder/norm/_0882_ ;
 wire \adder/norm/_0883_ ;
 wire net67;
 wire \adder/norm/_0885_ ;
 wire \adder/norm/_0886_ ;
 wire \adder/norm/_0887_ ;
 wire \adder/norm/_0888_ ;
 wire \adder/norm/_0889_ ;
 wire net66;
 wire \adder/norm/_0891_ ;
 wire \adder/norm/_0892_ ;
 wire net65;
 wire net64;
 wire \adder/norm/_0895_ ;
 wire \adder/norm/_0896_ ;
 wire \adder/norm/_0897_ ;
 wire \adder/norm/_0898_ ;
 wire \adder/norm/_0899_ ;
 wire \adder/norm/_0900_ ;
 wire \adder/norm/_0901_ ;
 wire \adder/norm/_0902_ ;
 wire \adder/norm/_0903_ ;
 wire \adder/norm/_0904_ ;
 wire \adder/norm/_0905_ ;
 wire \adder/norm/_0906_ ;
 wire net63;
 wire \adder/norm/_0908_ ;
 wire \adder/norm/_0909_ ;
 wire \adder/norm/_0910_ ;
 wire \adder/norm/_0911_ ;
 wire \adder/norm/_0912_ ;
 wire \adder/norm/_0913_ ;
 wire \adder/norm/_0914_ ;
 wire \adder/norm/_0915_ ;
 wire \adder/norm/_0916_ ;
 wire \adder/norm/_0917_ ;
 wire \adder/norm/_0918_ ;
 wire \adder/norm/_0919_ ;
 wire \adder/norm/_0920_ ;
 wire \adder/norm/_0921_ ;
 wire \adder/norm/_0922_ ;
 wire \adder/norm/_0923_ ;
 wire \adder/norm/_0924_ ;
 wire \adder/norm/_0925_ ;
 wire \adder/norm/_0926_ ;
 wire \adder/norm/_0927_ ;
 wire \adder/norm/_0928_ ;
 wire \adder/norm/_0929_ ;
 wire \adder/norm/_0930_ ;
 wire \adder/norm/_0931_ ;
 wire \adder/norm/_0932_ ;
 wire \adder/norm/_0933_ ;
 wire \adder/norm/_0934_ ;
 wire \adder/norm/_0935_ ;
 wire \adder/norm/_0936_ ;
 wire \adder/norm/_0937_ ;
 wire \adder/norm/_0938_ ;
 wire \adder/norm/_0939_ ;
 wire \adder/norm/_0940_ ;
 wire \adder/norm/_0941_ ;
 wire \adder/norm/_0942_ ;
 wire \adder/norm/_0943_ ;
 wire \adder/norm/_0944_ ;
 wire \adder/norm/_0945_ ;
 wire \adder/norm/_0946_ ;
 wire \adder/norm/_0947_ ;
 wire \adder/norm/_0948_ ;
 wire \adder/norm/_0949_ ;
 wire \adder/norm/_0950_ ;
 wire \adder/norm/_0951_ ;
 wire \adder/norm/_0952_ ;
 wire \adder/norm/_0953_ ;
 wire \adder/norm/_0954_ ;
 wire \adder/norm/_0955_ ;
 wire \adder/norm/_0956_ ;
 wire \adder/norm/_0957_ ;
 wire \adder/norm/_0958_ ;
 wire \adder/norm/_0959_ ;
 wire \adder/norm/_0960_ ;
 wire \adder/norm/_0961_ ;
 wire \adder/norm/_0962_ ;
 wire \adder/norm/_0963_ ;
 wire \adder/norm/_0964_ ;
 wire \adder/norm/_0965_ ;
 wire \adder/norm/_0966_ ;
 wire \adder/norm/_0967_ ;
 wire \adder/norm/_0968_ ;
 wire \adder/norm/_0969_ ;
 wire \adder/norm/_0970_ ;
 wire \adder/norm/_0971_ ;
 wire \adder/norm/_0972_ ;
 wire \adder/norm/_0973_ ;
 wire \adder/norm/_0974_ ;
 wire \adder/norm/_0975_ ;
 wire \adder/norm/_0976_ ;
 wire \adder/norm/_0977_ ;
 wire \adder/norm/_0978_ ;
 wire \adder/norm/_0979_ ;
 wire \adder/norm/_0980_ ;
 wire \adder/norm/_0981_ ;
 wire \adder/norm/_0982_ ;
 wire \adder/norm/_0983_ ;
 wire \adder/norm/_0984_ ;
 wire \adder/norm/_0985_ ;
 wire \adder/norm/_0986_ ;
 wire net62;
 wire net61;
 wire \adder/norm/_0989_ ;
 wire \adder/norm/_0990_ ;
 wire \adder/norm/_0991_ ;
 wire \adder/norm/_0992_ ;
 wire \adder/norm/_0993_ ;
 wire \adder/norm/_0994_ ;
 wire \adder/norm/_0995_ ;
 wire \adder/norm/_0996_ ;
 wire \adder/norm/_0997_ ;
 wire \adder/norm/_0998_ ;
 wire \adder/norm/_0999_ ;
 wire \adder/norm/_1000_ ;
 wire \adder/norm/_1001_ ;
 wire \adder/norm/_1002_ ;
 wire net60;
 wire net59;
 wire \adder/norm/_1005_ ;
 wire \adder/norm/_1006_ ;
 wire \adder/norm/_1007_ ;
 wire \adder/norm/_1008_ ;
 wire \adder/norm/_1009_ ;
 wire \adder/norm/_1010_ ;
 wire \adder/norm/_1011_ ;
 wire \adder/norm/_1012_ ;
 wire \adder/norm/_1013_ ;
 wire \adder/norm/_1014_ ;
 wire \adder/norm/_1015_ ;
 wire \adder/norm/_1016_ ;
 wire \adder/norm/_1017_ ;
 wire \adder/norm/_1018_ ;
 wire net58;
 wire \adder/norm/_1020_ ;
 wire \adder/norm/_1021_ ;
 wire \adder/norm/_1022_ ;
 wire \adder/norm/_1023_ ;
 wire \adder/norm/_1024_ ;
 wire \adder/norm/_1025_ ;
 wire \adder/norm/_1026_ ;
 wire \adder/norm/_1027_ ;
 wire \adder/norm/_1028_ ;
 wire \adder/norm/_1029_ ;
 wire \adder/norm/_1030_ ;
 wire \adder/norm/_1031_ ;
 wire \adder/norm/_1032_ ;
 wire \adder/norm/_1033_ ;
 wire \adder/norm/_1034_ ;
 wire \adder/norm/_1035_ ;
 wire \adder/norm/_1036_ ;
 wire \adder/norm/_1037_ ;
 wire \adder/norm/_1038_ ;
 wire \adder/norm/_1039_ ;
 wire \adder/norm/_1040_ ;
 wire \adder/norm/_1041_ ;
 wire \adder/norm/_1042_ ;
 wire \adder/norm/_1043_ ;
 wire \adder/norm/_1044_ ;
 wire \adder/norm/_1045_ ;
 wire \adder/norm/_1046_ ;
 wire \adder/norm/_1047_ ;
 wire \adder/norm/_1048_ ;
 wire \adder/norm/_1049_ ;
 wire \adder/norm/_1050_ ;
 wire \adder/norm/_1051_ ;
 wire \adder/norm/_1052_ ;
 wire \adder/norm/_1053_ ;
 wire \adder/norm/_1054_ ;
 wire \adder/norm/_1055_ ;
 wire \adder/norm/_1056_ ;
 wire \adder/norm/_1057_ ;
 wire \adder/norm/_1058_ ;
 wire \adder/norm/_1059_ ;
 wire \adder/norm/_1060_ ;
 wire \adder/norm/_1061_ ;
 wire \adder/norm/_1062_ ;
 wire \adder/norm/_1063_ ;
 wire \adder/norm/_1064_ ;
 wire \adder/norm/_1065_ ;
 wire \adder/norm/_1066_ ;
 wire \adder/norm/_1067_ ;
 wire \adder/norm/_1068_ ;
 wire net57;
 wire \adder/norm/_1070_ ;
 wire \adder/norm/_1071_ ;
 wire \adder/norm/_1072_ ;
 wire \adder/norm/_1073_ ;
 wire \adder/norm/_1074_ ;
 wire \adder/norm/_1075_ ;
 wire \adder/norm/_1076_ ;
 wire \adder/norm/_1077_ ;
 wire \adder/norm/_1078_ ;
 wire \adder/norm/_1079_ ;
 wire \adder/norm/_1080_ ;
 wire \adder/norm/_1081_ ;
 wire \adder/norm/_1082_ ;
 wire \adder/norm/_1083_ ;
 wire \adder/norm/_1084_ ;
 wire \adder/norm/_1085_ ;
 wire \adder/norm/_1086_ ;
 wire \adder/norm/_1087_ ;
 wire \adder/norm/_1088_ ;
 wire \adder/norm/_1089_ ;
 wire \adder/norm/_1090_ ;
 wire \adder/norm/_1091_ ;
 wire \adder/norm/_1092_ ;
 wire \adder/norm/_1093_ ;
 wire \adder/norm/_1094_ ;
 wire \adder/norm/_1095_ ;
 wire \adder/norm/_1096_ ;
 wire net56;
 wire \adder/norm/_1098_ ;
 wire \adder/norm/_1099_ ;
 wire \adder/norm/_1100_ ;
 wire \adder/norm/_1101_ ;
 wire \adder/norm/_1102_ ;
 wire \adder/norm/_1103_ ;
 wire \adder/norm/_1104_ ;
 wire \adder/norm/_1105_ ;
 wire \adder/norm/_1106_ ;
 wire \adder/norm/_1107_ ;
 wire \adder/norm/_1108_ ;
 wire \adder/norm/_1109_ ;
 wire \adder/norm/_1110_ ;
 wire \adder/norm/_1111_ ;
 wire \adder/norm/_1112_ ;
 wire \adder/norm/_1113_ ;
 wire \adder/norm/_1114_ ;
 wire \adder/norm/_1115_ ;
 wire \adder/norm/_1116_ ;
 wire \adder/norm/_1117_ ;
 wire \adder/norm/_1118_ ;
 wire \adder/norm/_1119_ ;
 wire \adder/norm/_1120_ ;
 wire \adder/norm/_1121_ ;
 wire \adder/norm/_1122_ ;
 wire \adder/norm/_1123_ ;
 wire \adder/norm/_1124_ ;
 wire \adder/norm/_1125_ ;
 wire \adder/norm/_1126_ ;
 wire \adder/norm/_1127_ ;
 wire \adder/norm/_1128_ ;
 wire \adder/norm/_1129_ ;
 wire \adder/norm/_1130_ ;
 wire \adder/norm/_1131_ ;
 wire \adder/norm/_1132_ ;
 wire \adder/norm/_1133_ ;
 wire \adder/norm/_1134_ ;
 wire \adder/norm/_1135_ ;
 wire \adder/norm/_1136_ ;
 wire \adder/norm/_1137_ ;
 wire \adder/norm/_1138_ ;
 wire \adder/norm/_1139_ ;
 wire \adder/norm/_1140_ ;
 wire \adder/norm/_1141_ ;
 wire \adder/norm/_1142_ ;
 wire \adder/norm/_1143_ ;
 wire \adder/norm/_1144_ ;
 wire \adder/norm/_1145_ ;
 wire \adder/norm/_1146_ ;
 wire \adder/norm/_1147_ ;
 wire \adder/norm/_1148_ ;
 wire \adder/norm/_1149_ ;
 wire \adder/norm/_1150_ ;
 wire \adder/norm/_1151_ ;
 wire \adder/norm/_1152_ ;
 wire \adder/norm/_1153_ ;
 wire \adder/norm/_1154_ ;
 wire \adder/norm/_1155_ ;
 wire \adder/norm/_1156_ ;
 wire \adder/norm/_1157_ ;
 wire \adder/norm/_1158_ ;
 wire \adder/norm/_1159_ ;
 wire \adder/norm/_1160_ ;
 wire \adder/norm/_1161_ ;
 wire \adder/norm/_1162_ ;
 wire \adder/norm/_1163_ ;
 wire \adder/norm/_1164_ ;
 wire \adder/norm/_1165_ ;
 wire \adder/norm/_1166_ ;
 wire \adder/norm/_1167_ ;
 wire \adder/norm/_1168_ ;
 wire \adder/norm/_1169_ ;
 wire \adder/norm/_1170_ ;
 wire \adder/norm/_1171_ ;
 wire \adder/norm/_1172_ ;
 wire \adder/norm/_1173_ ;
 wire \adder/norm/_1174_ ;
 wire \adder/norm/_1175_ ;
 wire \adder/norm/_1176_ ;
 wire \adder/norm/_1177_ ;
 wire \adder/norm/_1178_ ;
 wire \adder/norm/_1179_ ;
 wire \adder/norm/_1180_ ;
 wire \adder/norm/_1181_ ;
 wire net55;
 wire \adder/norm/_1183_ ;
 wire \adder/norm/_1184_ ;
 wire \adder/norm/_1185_ ;
 wire \adder/norm/_1186_ ;
 wire \adder/norm/_1187_ ;
 wire \adder/norm/_1188_ ;
 wire \adder/norm/_1189_ ;
 wire \adder/norm/_1190_ ;
 wire \adder/norm/_1191_ ;
 wire \adder/norm/_1192_ ;
 wire \adder/norm/_1193_ ;
 wire \adder/norm/_1194_ ;
 wire \adder/norm/_1195_ ;
 wire \adder/norm/_1196_ ;
 wire \adder/norm/_1197_ ;
 wire \adder/norm/_1198_ ;
 wire \adder/norm/_1199_ ;
 wire \adder/norm/_1200_ ;
 wire \adder/norm/_1201_ ;
 wire \adder/norm/_1202_ ;
 wire \adder/norm/_1203_ ;
 wire \adder/norm/_1204_ ;
 wire \adder/norm/_1205_ ;
 wire \adder/norm/_1206_ ;
 wire \adder/norm/_1207_ ;
 wire \adder/norm/_1208_ ;
 wire \adder/norm/_1209_ ;
 wire \adder/norm/_1210_ ;
 wire \adder/norm/_1211_ ;
 wire \adder/norm/_1212_ ;
 wire \adder/norm/_1213_ ;
 wire \adder/norm/_1214_ ;
 wire \adder/norm/_1215_ ;
 wire \adder/norm/_1216_ ;
 wire \adder/norm/_1217_ ;
 wire \adder/norm/_1218_ ;
 wire \adder/norm/_1219_ ;
 wire \adder/norm/_1220_ ;
 wire \adder/norm/_1221_ ;
 wire \adder/norm/_1222_ ;
 wire \adder/norm/_1223_ ;
 wire \adder/norm/_1224_ ;
 wire \adder/norm/_1225_ ;
 wire \adder/norm/_1226_ ;
 wire \adder/norm/_1227_ ;
 wire \adder/norm/_1228_ ;
 wire \adder/norm/_1229_ ;
 wire \adder/norm/_1230_ ;
 wire \adder/norm/_1231_ ;
 wire net54;
 wire \adder/norm/_1233_ ;
 wire \adder/norm/_1234_ ;
 wire \adder/norm/_1235_ ;
 wire \adder/norm/_1236_ ;
 wire \adder/norm/_1237_ ;
 wire \adder/norm/_1238_ ;
 wire \adder/norm/_1239_ ;
 wire \adder/norm/_1240_ ;
 wire \adder/norm/_1241_ ;
 wire \adder/norm/_1242_ ;
 wire \adder/norm/_1243_ ;
 wire \adder/norm/_1244_ ;
 wire \adder/norm/_1245_ ;
 wire \adder/norm/_1246_ ;
 wire \adder/norm/_1247_ ;
 wire \adder/norm/_1248_ ;
 wire \adder/norm/_1249_ ;
 wire \adder/norm/_1250_ ;
 wire \adder/norm/_1251_ ;
 wire \adder/norm/_1252_ ;
 wire \adder/norm/_1253_ ;
 wire \adder/norm/_1254_ ;
 wire \adder/norm/_1255_ ;
 wire \adder/norm/_1256_ ;
 wire \adder/norm/_1257_ ;
 wire \adder/norm/_1258_ ;
 wire \adder/norm/_1259_ ;
 wire \adder/norm/_1260_ ;
 wire \adder/norm/_1261_ ;
 wire \adder/norm/_1262_ ;
 wire \adder/norm/_1263_ ;
 wire \adder/norm/_1264_ ;
 wire \adder/norm/_1265_ ;
 wire \adder/norm/_1266_ ;
 wire \adder/norm/_1267_ ;
 wire \adder/norm/_1268_ ;
 wire \adder/norm/_1269_ ;
 wire \adder/norm/_1270_ ;
 wire \adder/norm/_1271_ ;
 wire \adder/norm/_1272_ ;
 wire \adder/norm/_1273_ ;
 wire net53;
 wire \adder/norm/_1275_ ;
 wire \adder/norm/_1276_ ;
 wire \adder/norm/_1277_ ;
 wire \adder/norm/_1278_ ;
 wire \adder/norm/_1279_ ;
 wire \adder/norm/_1280_ ;
 wire \adder/norm/_1281_ ;
 wire \adder/norm/_1282_ ;
 wire \adder/norm/_1283_ ;
 wire \adder/norm/_1284_ ;
 wire \adder/norm/_1285_ ;
 wire \adder/norm/_1286_ ;
 wire \adder/norm/_1287_ ;
 wire \adder/norm/_1288_ ;
 wire \adder/norm/_1289_ ;
 wire \adder/norm/_1290_ ;
 wire \adder/norm/_1291_ ;
 wire \adder/norm/_1292_ ;
 wire \adder/norm/_1293_ ;
 wire \adder/norm/_1294_ ;
 wire \adder/norm/_1295_ ;
 wire \adder/norm/_1296_ ;
 wire \adder/norm/_1297_ ;
 wire \adder/norm/_1298_ ;
 wire \adder/norm/_1299_ ;
 wire \adder/norm/_1300_ ;
 wire \adder/norm/_1301_ ;
 wire \adder/norm/_1302_ ;
 wire \adder/norm/_1303_ ;
 wire \adder/norm/_1304_ ;
 wire \adder/norm/_1305_ ;
 wire \adder/norm/_1306_ ;
 wire \adder/norm/_1307_ ;
 wire \adder/norm/_1308_ ;
 wire \adder/norm/_1309_ ;
 wire \adder/norm/_1310_ ;
 wire \adder/norm/_1311_ ;
 wire \adder/norm/_1312_ ;
 wire \adder/norm/_1313_ ;
 wire \adder/norm/_1314_ ;
 wire \adder/norm/_1315_ ;
 wire \adder/norm/_1316_ ;
 wire \adder/norm/_1317_ ;
 wire \adder/norm/_1318_ ;
 wire \adder/norm/_1319_ ;
 wire \adder/norm/_1320_ ;
 wire \adder/norm/_1321_ ;
 wire \adder/norm/_1322_ ;
 wire \adder/norm/_1323_ ;
 wire \adder/norm/_1324_ ;
 wire \adder/norm/_1325_ ;
 wire \adder/norm/_1326_ ;
 wire \adder/norm/_1327_ ;
 wire \adder/norm/_1328_ ;
 wire \adder/norm/_1329_ ;
 wire \adder/norm/_1330_ ;
 wire \adder/norm/_1331_ ;
 wire \adder/norm/_1332_ ;
 wire \adder/norm/_1333_ ;
 wire \adder/norm/_1334_ ;
 wire \adder/norm/_1335_ ;
 wire \adder/norm/_1336_ ;
 wire \adder/norm/_1337_ ;
 wire \adder/norm/_1338_ ;
 wire \adder/norm/_1339_ ;
 wire \adder/norm/_1340_ ;
 wire \adder/norm/_1341_ ;
 wire \adder/norm/_1342_ ;
 wire \adder/norm/_1343_ ;
 wire \adder/norm/_1344_ ;
 wire \adder/norm/_1345_ ;
 wire \adder/norm/_1346_ ;
 wire \adder/norm/_1347_ ;
 wire \adder/norm/_1348_ ;
 wire \adder/norm/_1349_ ;
 wire \adder/norm/_1350_ ;
 wire \adder/norm/_1351_ ;
 wire \adder/norm/_1352_ ;
 wire \adder/norm/_1353_ ;
 wire \adder/norm/_1354_ ;
 wire \adder/norm/_1355_ ;
 wire \adder/norm/_1356_ ;
 wire \adder/norm/_1357_ ;
 wire \adder/norm/_1358_ ;
 wire \adder/norm/_1359_ ;
 wire \adder/norm/_1360_ ;
 wire \adder/norm/_1361_ ;
 wire \adder/norm/_1362_ ;
 wire \adder/norm/_1363_ ;
 wire \adder/norm/_1364_ ;
 wire \adder/norm/_1365_ ;
 wire \adder/norm/_1366_ ;
 wire \adder/norm/_1367_ ;
 wire \adder/norm/_1368_ ;
 wire \adder/norm/_1369_ ;
 wire \adder/norm/_1370_ ;
 wire \adder/norm/_1371_ ;
 wire \adder/norm/_1372_ ;
 wire \adder/norm/_1373_ ;
 wire \adder/norm/_1374_ ;
 wire \adder/norm/_1375_ ;
 wire \adder/norm/_1376_ ;
 wire \adder/norm/_1377_ ;
 wire \adder/norm/_1378_ ;
 wire \adder/norm/_1379_ ;
 wire \adder/norm/_1380_ ;
 wire \adder/norm/_1381_ ;
 wire \adder/norm/_1382_ ;
 wire \adder/norm/_1383_ ;
 wire \adder/norm/_1384_ ;
 wire \adder/norm/_1385_ ;
 wire \adder/norm/_1386_ ;
 wire \adder/norm/_1387_ ;
 wire \adder/norm/_1388_ ;
 wire \adder/norm/_1389_ ;
 wire \adder/norm/_1390_ ;
 wire \adder/norm/_1391_ ;
 wire \adder/norm/_1392_ ;
 wire \adder/norm/_1393_ ;
 wire \adder/norm/_1394_ ;
 wire \adder/norm/_1395_ ;
 wire \adder/norm/_1396_ ;
 wire \adder/norm/_1397_ ;
 wire \adder/norm/_1398_ ;
 wire \adder/norm/_1399_ ;
 wire \adder/norm/_1400_ ;
 wire \adder/norm/_1401_ ;
 wire \adder/norm/_1402_ ;
 wire \adder/norm/_1403_ ;
 wire \adder/norm/_1404_ ;
 wire \adder/norm/_1405_ ;
 wire \adder/norm/_1406_ ;
 wire \adder/norm/_1407_ ;
 wire \adder/norm/_1408_ ;
 wire \adder/norm/_1409_ ;
 wire \adder/norm/_1410_ ;
 wire \adder/norm/_1411_ ;
 wire \adder/norm/_1412_ ;
 wire \adder/norm/_1413_ ;
 wire \adder/norm/_1414_ ;
 wire \adder/norm/_1415_ ;
 wire \adder/norm/_1416_ ;
 wire \adder/norm/_1417_ ;
 wire \adder/norm/_1418_ ;
 wire \adder/norm/_1419_ ;
 wire \adder/norm/_1420_ ;
 wire \adder/norm/_1421_ ;
 wire \adder/norm/_1422_ ;
 wire \adder/norm/_1423_ ;
 wire \adder/norm/_1424_ ;
 wire \adder/norm/_1425_ ;
 wire \adder/norm/_1426_ ;
 wire \adder/norm/_1427_ ;
 wire \adder/norm/_1428_ ;
 wire \adder/norm/_1429_ ;
 wire \adder/norm/_1430_ ;
 wire \adder/norm/_1431_ ;
 wire \adder/norm/_1432_ ;
 wire \adder/norm/_1433_ ;
 wire \adder/norm/_1434_ ;
 wire \adder/norm/_1435_ ;
 wire \adder/norm/_1436_ ;
 wire \adder/norm/_1437_ ;
 wire \adder/norm/_1438_ ;
 wire \adder/norm/_1439_ ;
 wire \adder/norm/_1440_ ;
 wire \adder/norm/_1441_ ;
 wire \adder/norm/_1442_ ;
 wire \adder/norm/_1443_ ;
 wire \adder/norm/_1444_ ;
 wire net52;
 wire \adder/norm/_1446_ ;
 wire \adder/norm/_1447_ ;
 wire \adder/norm/_1448_ ;
 wire \adder/norm/_1449_ ;
 wire \adder/norm/_1450_ ;
 wire \adder/norm/_1451_ ;
 wire \adder/norm/_1452_ ;
 wire \adder/norm/_1453_ ;
 wire \adder/norm/_1454_ ;
 wire \adder/norm/_1455_ ;
 wire \adder/norm/_1456_ ;
 wire \adder/norm/_1457_ ;
 wire \adder/norm/_1458_ ;
 wire \adder/norm/_1459_ ;
 wire \adder/norm/_1460_ ;
 wire \adder/norm/_1461_ ;
 wire \adder/norm/_1462_ ;
 wire \adder/norm/_1463_ ;
 wire \adder/norm/_1464_ ;
 wire \adder/norm/_1465_ ;
 wire \adder/norm/_1466_ ;
 wire \adder/norm/_1467_ ;
 wire \adder/norm/_1468_ ;
 wire \adder/norm/_1469_ ;
 wire \adder/norm/_1470_ ;
 wire \adder/norm/_1471_ ;
 wire \adder/norm/_1472_ ;
 wire \adder/norm/_1473_ ;
 wire \adder/norm/_1474_ ;
 wire \adder/norm/_1475_ ;
 wire \adder/norm/LOD/_000_ ;
 wire \adder/norm/LOD/_001_ ;
 wire \adder/norm/LOD/_002_ ;
 wire \adder/norm/LOD/_003_ ;
 wire \adder/norm/LOD/_004_ ;
 wire \adder/norm/LOD/_005_ ;
 wire \adder/norm/LOD/_006_ ;
 wire \adder/norm/LOD/_007_ ;
 wire \adder/norm/LOD/_008_ ;
 wire \adder/norm/LOD/_009_ ;
 wire \adder/norm/LOD/_010_ ;
 wire \adder/norm/LOD/_011_ ;
 wire \adder/norm/LOD/_012_ ;
 wire \adder/norm/LOD/_013_ ;
 wire \adder/norm/LOD/_014_ ;
 wire \adder/norm/LOD/_015_ ;
 wire \adder/norm/LOD/_016_ ;
 wire \adder/norm/LOD/_017_ ;
 wire \adder/norm/LOD/_018_ ;
 wire \adder/norm/LOD/_019_ ;
 wire \adder/norm/LOD/_020_ ;
 wire \adder/norm/LOD/_021_ ;
 wire \adder/norm/LOD/_022_ ;
 wire \adder/norm/LOD/_023_ ;
 wire \adder/norm/LOD/_024_ ;
 wire \adder/norm/LOD/_025_ ;
 wire \adder/norm/LOD/_026_ ;
 wire \adder/norm/LOD/_027_ ;
 wire \adder/norm/LOD/_028_ ;
 wire \adder/norm/LOD/_029_ ;
 wire \adder/norm/LOD/_030_ ;
 wire \adder/norm/LOD/_031_ ;
 wire \adder/norm/LOD/_032_ ;
 wire \adder/norm/LOD/_033_ ;
 wire \adder/norm/LOD/_034_ ;
 wire \adder/norm/LOD/_035_ ;
 wire \adder/norm/LOD/_036_ ;
 wire \adder/norm/LOD/_037_ ;
 wire \adder/norm/LOD/_038_ ;
 wire \adder/norm/LOD/_039_ ;
 wire \adder/norm/LOD/_040_ ;
 wire \adder/norm/LOD/_041_ ;
 wire \adder/norm/LOD/_042_ ;
 wire \adder/norm/LOD/_043_ ;
 wire \adder/norm/LOD/_044_ ;
 wire \adder/norm/LOD/_045_ ;
 wire \adder/norm/LOD/_046_ ;
 wire \adder/norm/LOD/_047_ ;
 wire \adder/norm/LOD/_048_ ;
 wire \adder/norm/LOD/_049_ ;
 wire \adder/norm/LOD/_050_ ;
 wire \adder/norm/LOD/_051_ ;
 wire \adder/norm/LOD/_052_ ;
 wire \adder/norm/LOD/_053_ ;
 wire \adder/norm/LOD/_054_ ;
 wire \adder/norm/LOD/_055_ ;
 wire \adder/norm/LOD/_056_ ;
 wire \adder/norm/LOD/_057_ ;
 wire \adder/norm/LOD/_058_ ;
 wire \adder/norm/LOD/_059_ ;
 wire \adder/norm/LOD/_060_ ;
 wire \adder/norm/LOD/_061_ ;
 wire \adder/norm/LOD/_062_ ;
 wire \adder/norm/LOD/_063_ ;
 wire \adder/norm/LOD/_064_ ;
 wire \adder/norm/LOD/_065_ ;
 wire \adder/norm/LOD/_066_ ;
 wire \adder/norm/LOD/_067_ ;
 wire \adder/norm/LOD/_068_ ;
 wire \adder/norm/LOD/_069_ ;
 wire \adder/norm/LOD/_070_ ;
 wire \adder/norm/LOD/_071_ ;
 wire \adder/norm/LOD/_072_ ;
 wire \adder/norm/LOD/_073_ ;
 wire \adder/norm/LOD/_074_ ;
 wire \adder/norm/LOD/_075_ ;
 wire \adder/norm/LOD/_076_ ;
 wire \adder/norm/LOD/_077_ ;
 wire \adder/norm/LOD/_078_ ;
 wire \adder/norm/LOD/_079_ ;
 wire \adder/norm/LOD/_080_ ;
 wire \adder/norm/LOD/_081_ ;
 wire \adder/norm/LOD/_082_ ;
 wire \adder/norm/LOD/_083_ ;
 wire \adder/norm/LOD/_084_ ;
 wire \adder/norm/LOD/_085_ ;
 wire \adder/norm/LOD/_086_ ;
 wire \adder/norm/LOD/_087_ ;
 wire \adder/norm/LOD/_088_ ;
 wire \adder/norm/LOD/_089_ ;
 wire \adder/norm/LOD/_090_ ;
 wire \adder/norm/LOD/_091_ ;
 wire \adder/norm/LOD/_092_ ;
 wire \adder/norm/LOD/_093_ ;
 wire \adder/norm/LOD/_094_ ;
 wire \adder/norm/LOD/_095_ ;
 wire \adder/norm/LOD/_096_ ;
 wire \adder/norm/LOD/_097_ ;
 wire \adder/norm/LOD/_098_ ;
 wire \adder/norm/LOD/_099_ ;
 wire \adder/norm/LOD/_100_ ;
 wire \adder/norm/LOD/_101_ ;
 wire \adder/norm/LOD/_102_ ;
 wire \adder/norm/LOD/_103_ ;
 wire \adder/norm/LOD/_104_ ;
 wire \adder/norm/LOD/_105_ ;
 wire \adder/norm/LOD/_106_ ;
 wire \adder/norm/LOD/_107_ ;
 wire \adder/norm/LOD/_108_ ;
 wire \adder/norm/LOD/_109_ ;
 wire \adder/norm/LOD/_110_ ;
 wire \adder/norm/LOD/_111_ ;
 wire \adder/norm/LOD/_112_ ;
 wire \adder/norm/LOD/_113_ ;
 wire \adder/norm/LOD/_114_ ;
 wire \adder/norm/LOD/_115_ ;
 wire \adder/norm/LOD/_116_ ;
 wire \adder/norm/LOD/_117_ ;
 wire \adder/norm/LOD/_118_ ;
 wire \adder/norm/LOD/_119_ ;
 wire \adder/norm/LOD/_120_ ;
 wire \adder/norm/LOD/_121_ ;
 wire \adder/norm/LOD/_122_ ;
 wire \adder/norm/LOD/_123_ ;
 wire \adder/norm/LOD/_124_ ;
 wire \adder/norm/LOD/_125_ ;
 wire \adder/norm/LOD/_126_ ;
 wire \adder/norm/LOD/_127_ ;
 wire \adder/norm/LOD/_128_ ;
 wire \adder/norm/LOD/_129_ ;
 wire \adder/norm/LOD/_130_ ;
 wire \adder/norm/LOD/_131_ ;
 wire \adder/norm/LOD/_132_ ;
 wire \adder/norm/LOD/_133_ ;
 wire \adder/norm/LOD/_134_ ;
 wire \adder/norm/LOD/_135_ ;
 wire \adder/norm/LOD/_136_ ;
 wire \adder/norm/LOD/_137_ ;
 wire \adder/norm/LOD/_138_ ;
 wire \adder/norm/LOD/_139_ ;
 wire \adder/norm/LOD/_140_ ;
 wire \adder/norm/LOD/_141_ ;
 wire \adder/norm/LOD/_142_ ;
 wire \adder/norm/LOD/_143_ ;
 wire \adder/norm/LOD/_144_ ;
 wire \adder/norm/LOD/_145_ ;
 wire \adder/norm/LOD/_146_ ;
 wire \adder/norm/LOD/_147_ ;
 wire \adder/norm/LOD/_148_ ;
 wire \adder/norm/LOD/_149_ ;
 wire \adder/norm/LOD/_150_ ;
 wire \adder/norm/LOD/_151_ ;
 wire \adder/norm/LOD/_152_ ;
 wire \adder/norm/LOD/_153_ ;
 wire \adder/norm/LOD/_154_ ;
 wire \adder/norm/LOD/_155_ ;
 wire \adder/norm/LOD/_156_ ;
 wire \converter/_000_ ;
 wire \converter/_001_ ;
 wire \converter/_002_ ;
 wire \converter/_003_ ;
 wire \converter/_004_ ;
 wire \converter/_005_ ;
 wire \converter/_006_ ;
 wire \converter/_007_ ;
 wire \converter/_008_ ;
 wire \converter/_009_ ;
 wire \converter/_010_ ;
 wire \converter/_011_ ;
 wire \converter/_012_ ;
 wire \converter/_013_ ;
 wire \converter/_014_ ;
 wire \converter/_015_ ;
 wire \converter/_016_ ;
 wire \converter/_017_ ;
 wire \converter/_018_ ;
 wire \converter/_019_ ;
 wire \converter/_020_ ;
 wire \converter/_021_ ;
 wire \converter/_022_ ;
 wire \converter/_023_ ;
 wire \converter/_024_ ;
 wire \converter/_025_ ;
 wire \converter/_026_ ;
 wire \converter/_027_ ;
 wire \converter/_028_ ;
 wire \converter/_029_ ;
 wire \converter/_030_ ;
 wire \converter/_031_ ;
 wire \converter/_032_ ;
 wire \converter/_033_ ;
 wire \converter/_034_ ;
 wire \converter/_035_ ;
 wire \converter/_036_ ;
 wire \converter/_037_ ;
 wire \converter/_038_ ;
 wire \converter/_039_ ;
 wire \converter/_040_ ;
 wire \converter/_041_ ;
 wire \converter/_042_ ;
 wire \converter/_043_ ;
 wire \converter/_044_ ;
 wire \converter/_045_ ;
 wire \converter/_046_ ;
 wire \converter/_047_ ;
 wire \converter/_048_ ;
 wire \converter/_049_ ;
 wire \converter/_050_ ;
 wire \converter/_051_ ;
 wire \converter/_052_ ;
 wire \converter/_053_ ;
 wire \converter/_054_ ;
 wire \converter/_055_ ;
 wire \converter/_056_ ;
 wire \converter/_057_ ;
 wire \converter/_058_ ;
 wire \converter/_059_ ;
 wire \converter/_060_ ;
 wire \converter/_061_ ;
 wire \converter/_062_ ;
 wire \converter/_063_ ;
 wire \converter/_064_ ;
 wire \converter/_065_ ;
 wire \converter/_066_ ;
 wire \converter/_067_ ;
 wire \converter/_068_ ;
 wire \converter/_069_ ;
 wire \converter/_070_ ;
 wire \converter/_071_ ;
 wire \converter/_072_ ;
 wire \converter/_073_ ;
 wire \converter/_074_ ;
 wire \converter/_075_ ;
 wire \converter/_076_ ;
 wire \converter/_077_ ;
 wire \converter/_078_ ;
 wire \converter/_079_ ;
 wire \converter/_080_ ;
 wire \converter/_081_ ;
 wire \converter/_082_ ;
 wire \converter/_083_ ;
 wire \converter/_084_ ;
 wire \converter/_085_ ;
 wire \converter/_086_ ;
 wire \converter/_087_ ;
 wire \converter/_088_ ;
 wire \converter/_089_ ;
 wire \converter/_090_ ;
 wire \converter/_091_ ;
 wire \converter/_092_ ;
 wire \converter/_093_ ;
 wire \converter/_094_ ;
 wire \converter/_095_ ;
 wire \converter/_096_ ;
 wire \converter/_097_ ;
 wire net23;
 wire \converter/_099_ ;
 wire \converter/_100_ ;
 wire net22;
 wire net21;
 wire \converter/_103_ ;
 wire \converter/_104_ ;
 wire \converter/_105_ ;
 wire net20;
 wire \converter/_107_ ;
 wire \converter/_108_ ;
 wire \converter/_109_ ;
 wire \converter/_110_ ;
 wire \converter/_111_ ;
 wire \converter/_112_ ;
 wire net19;
 wire \converter/_114_ ;
 wire net18;
 wire \converter/_116_ ;
 wire \converter/_117_ ;
 wire \converter/_118_ ;
 wire \converter/_119_ ;
 wire \converter/_120_ ;
 wire \converter/_121_ ;
 wire \converter/_122_ ;
 wire \converter/_123_ ;
 wire \converter/_124_ ;
 wire \converter/_125_ ;
 wire \converter/_126_ ;
 wire \converter/_127_ ;
 wire \converter/_128_ ;
 wire \converter/_129_ ;
 wire \converter/_130_ ;
 wire \converter/_131_ ;
 wire \converter/_132_ ;
 wire \converter/_133_ ;
 wire \converter/_134_ ;
 wire \converter/_135_ ;
 wire \converter/_136_ ;
 wire \converter/_137_ ;
 wire \converter/_138_ ;
 wire \converter/_139_ ;
 wire \converter/_140_ ;
 wire \converter/_141_ ;
 wire \converter/_142_ ;
 wire \converter/_143_ ;
 wire \converter/_144_ ;
 wire \converter/_145_ ;
 wire net17;
 wire net16;
 wire \converter/_148_ ;
 wire \converter/_149_ ;
 wire \converter/_150_ ;
 wire net15;
 wire \converter/_152_ ;
 wire \converter/_153_ ;
 wire \converter/_154_ ;
 wire \converter/_155_ ;
 wire \converter/_156_ ;
 wire \converter/_157_ ;
 wire \converter/_158_ ;
 wire \converter/_159_ ;
 wire \converter/_160_ ;
 wire net239;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;

 NOR2_X1 \adder/_20_  (.A1(\operand_fp16_fp32[29] ),
    .A2(\operand_fp16_fp32[27] ),
    .ZN(\adder/_00_ ));
 NOR2_X1 \adder/_21_  (.A1(net6),
    .A2(\operand_fp16_fp32[29] ),
    .ZN(\adder/_01_ ));
 AND2_X1 \adder/_22_  (.A1(\adder/_00_ ),
    .A2(\adder/_01_ ),
    .ZN(\adder/_02_ ));
 INV_X1 \adder/_23_  (.A(\operand_fp16_fp32[24] ),
    .ZN(\adder/_03_ ));
 INV_X1 \adder/_24_  (.A(\operand_fp16_fp32[23] ),
    .ZN(\adder/_04_ ));
 NAND2_X1 \adder/_25_  (.A1(\adder/_03_ ),
    .A2(\adder/_04_ ),
    .ZN(\adder/_05_ ));
 INV_X1 \adder/_26_  (.A(\operand_fp16_fp32[26] ),
    .ZN(\adder/_06_ ));
 INV_X1 \adder/_27_  (.A(\operand_fp16_fp32[25] ),
    .ZN(\adder/_07_ ));
 NAND2_X1 \adder/_28_  (.A1(\adder/_06_ ),
    .A2(\adder/_07_ ),
    .ZN(\adder/_08_ ));
 NOR2_X1 \adder/_29_  (.A1(\adder/_05_ ),
    .A2(\adder/_08_ ),
    .ZN(\adder/_09_ ));
 NAND2_X1 \adder/_30_  (.A1(\adder/_02_ ),
    .A2(\adder/_09_ ),
    .ZN(\adder/hb_a_d ));
 NOR2_X1 \adder/_31_  (.A1(net37),
    .A2(net36),
    .ZN(\adder/_10_ ));
 NOR2_X1 \adder/_32_  (.A1(net40),
    .A2(net38),
    .ZN(\adder/_11_ ));
 AND2_X1 \adder/_33_  (.A1(\adder/_10_ ),
    .A2(\adder/_11_ ),
    .ZN(\adder/_12_ ));
 INV_X1 \adder/_34_  (.A(net33),
    .ZN(\adder/_13_ ));
 INV_X1 \adder/_35_  (.A(net32),
    .ZN(\adder/_14_ ));
 NAND2_X1 \adder/_36_  (.A1(\adder/_13_ ),
    .A2(\adder/_14_ ),
    .ZN(\adder/_15_ ));
 INV_X1 \adder/_37_  (.A(net35),
    .ZN(\adder/_16_ ));
 INV_X1 \adder/_38_  (.A(net34),
    .ZN(\adder/_17_ ));
 NAND2_X1 \adder/_39_  (.A1(\adder/_16_ ),
    .A2(\adder/_17_ ),
    .ZN(\adder/_18_ ));
 NOR2_X1 \adder/_40_  (.A1(\adder/_15_ ),
    .A2(\adder/_18_ ),
    .ZN(\adder/_19_ ));
 NAND2_X1 \adder/_41_  (.A1(\adder/_12_ ),
    .A2(\adder/_19_ ),
    .ZN(\adder/hb_b_d ));
 BUF_X16 max_cap85 (.A(\adder/adder/_0451_ ),
    .Z(net85));
 NOR2_X1 \adder/adder/_1108_  (.A1(\adder/adder/_0307_ ),
    .A2(\operand_fp16_fp32[21] ),
    .ZN(\adder/adder/_0308_ ));
 INV_X1 \adder/adder/_1109_  (.A(\operand_fp16_fp32[21] ),
    .ZN(\adder/adder/_0309_ ));
 NOR2_X1 \adder/adder/_1110_  (.A1(\adder/adder/_0309_ ),
    .A2(net30),
    .ZN(\adder/adder/_0310_ ));
 NOR2_X1 \adder/adder/_1111_  (.A1(\adder/adder/_0308_ ),
    .A2(\adder/adder/_0310_ ),
    .ZN(\adder/adder/_0311_ ));
 INV_X1 \adder/adder/_1112_  (.A(\adder/adder/_0311_ ),
    .ZN(\adder/adder/_0312_ ));
 INV_X1 \adder/adder/_1113_  (.A(\operand_fp16_fp32[20] ),
    .ZN(\adder/adder/_0313_ ));
 NOR2_X1 \adder/adder/_1114_  (.A1(\adder/adder/_0313_ ),
    .A2(net29),
    .ZN(\adder/adder/_0314_ ));
 INV_X1 \adder/adder/_1115_  (.A(net29),
    .ZN(\adder/adder/_0315_ ));
 NOR2_X1 \adder/adder/_1116_  (.A1(\adder/adder/_0315_ ),
    .A2(\operand_fp16_fp32[20] ),
    .ZN(\adder/adder/_0316_ ));
 NOR4_X1 \adder/adder/_1117_  (.A1(\adder/adder/_0306_ ),
    .A2(\adder/adder/_0312_ ),
    .A3(\adder/adder/_0314_ ),
    .A4(\adder/adder/_0316_ ),
    .ZN(\adder/adder/_0317_ ));
 INV_X1 \adder/adder/_1118_  (.A(\adder/adder/_0317_ ),
    .ZN(\adder/adder/_0318_ ));
 INV_X1 \adder/adder/_1119_  (.A(\operand_fp16_fp32[17] ),
    .ZN(\adder/adder/_0319_ ));
 BUF_X16 wire84 (.A(\adder/norm/_0670_ ),
    .Z(net84));
 XNOR2_X1 \adder/adder/_1121_  (.A(\adder/adder/_0319_ ),
    .B(net25),
    .ZN(\adder/adder/_0321_ ));
 INV_X1 \adder/adder/_1122_  (.A(net27),
    .ZN(\adder/adder/_0322_ ));
 OR2_X1 \adder/adder/_1123_  (.A1(\adder/adder/_0322_ ),
    .A2(\operand_fp16_fp32[19] ),
    .ZN(\adder/adder/_0323_ ));
 NAND2_X1 \adder/adder/_1124_  (.A1(\adder/adder/_0322_ ),
    .A2(\operand_fp16_fp32[19] ),
    .ZN(\adder/adder/_0324_ ));
 AND2_X1 \adder/adder/_1125_  (.A1(\adder/adder/_0323_ ),
    .A2(\adder/adder/_0324_ ),
    .ZN(\adder/adder/_0325_ ));
 INV_X1 \adder/adder/_1126_  (.A(net26),
    .ZN(\adder/adder/_0326_ ));
 NOR2_X1 \adder/adder/_1127_  (.A1(\adder/adder/_0326_ ),
    .A2(\operand_fp16_fp32[18] ),
    .ZN(\adder/adder/_0327_ ));
 INV_X1 \adder/adder/_1128_  (.A(\adder/adder/_0327_ ),
    .ZN(\adder/adder/_0328_ ));
 NAND2_X1 \adder/adder/_1129_  (.A1(\adder/adder/_0326_ ),
    .A2(\operand_fp16_fp32[18] ),
    .ZN(\adder/adder/_0329_ ));
 NAND3_X1 \adder/adder/_1130_  (.A1(\adder/adder/_0325_ ),
    .A2(\adder/adder/_0328_ ),
    .A3(\adder/adder/_0329_ ),
    .ZN(\adder/adder/_0330_ ));
 INV_X1 \adder/adder/_1131_  (.A(net24),
    .ZN(\adder/adder/_0331_ ));
 NAND2_X1 \adder/adder/_1132_  (.A1(\adder/adder/_0331_ ),
    .A2(\operand_fp16_fp32[16] ),
    .ZN(\adder/adder/_0332_ ));
 INV_X1 \adder/adder/_1133_  (.A(\operand_fp16_fp32[16] ),
    .ZN(\adder/adder/_0333_ ));
 NAND2_X1 \adder/adder/_1134_  (.A1(\adder/adder/_0333_ ),
    .A2(net24),
    .ZN(\adder/adder/_0334_ ));
 NAND2_X1 \adder/adder/_1135_  (.A1(\adder/adder/_0332_ ),
    .A2(\adder/adder/_0334_ ),
    .ZN(\adder/adder/_0335_ ));
 NOR4_X1 \adder/adder/_1136_  (.A1(\adder/adder/_0318_ ),
    .A2(\adder/adder/_0321_ ),
    .A3(\adder/adder/_0330_ ),
    .A4(\adder/adder/_0335_ ),
    .ZN(\adder/adder/_0336_ ));
 NAND2_X1 \adder/adder/_1137_  (.A1(\adder/adder/_0299_ ),
    .A2(\adder/adder/_0336_ ),
    .ZN(\adder/adder/_0337_ ));
 INV_X1 \adder/adder/_1138_  (.A(\adder/hb_b_d ),
    .ZN(\adder/adder/_0338_ ));
 NOR2_X1 \adder/adder/_1139_  (.A1(\adder/adder/_0338_ ),
    .A2(\adder/hb_a_d ),
    .ZN(\adder/adder/_0339_ ));
 AOI21_X1 \adder/adder/_1140_  (.A(\adder/adder/_0339_ ),
    .B1(\adder/adder/_0301_ ),
    .B2(\adder/adder/_0303_ ),
    .ZN(\adder/adder/_0340_ ));
 AOI21_X1 \adder/adder/_1141_  (.A(\adder/adder/_0308_ ),
    .B1(\adder/adder/_0311_ ),
    .B2(\adder/adder/_0316_ ),
    .ZN(\adder/adder/_0341_ ));
 INV_X1 \adder/adder/_1142_  (.A(\adder/adder/_0325_ ),
    .ZN(\adder/adder/_0342_ ));
 NOR2_X1 \adder/adder/_1143_  (.A1(\adder/adder/_0321_ ),
    .A2(\adder/adder/_0334_ ),
    .ZN(\adder/adder/_0343_ ));
 AOI21_X1 \adder/adder/_1144_  (.A(\adder/adder/_0343_ ),
    .B1(\adder/adder/_0319_ ),
    .B2(net25),
    .ZN(\adder/adder/_0344_ ));
 OAI221_X1 \adder/adder/_1145_  (.A(\adder/adder/_0323_ ),
    .B1(\adder/adder/_0342_ ),
    .B2(\adder/adder/_0328_ ),
    .C1(\adder/adder/_0344_ ),
    .C2(\adder/adder/_0330_ ),
    .ZN(\adder/adder/_0345_ ));
 INV_X1 \adder/adder/_1146_  (.A(\adder/adder/_0345_ ),
    .ZN(\adder/adder/_0346_ ));
 OAI221_X1 \adder/adder/_1147_  (.A(\adder/adder/_0340_ ),
    .B1(\adder/adder/_0306_ ),
    .B2(\adder/adder/_0341_ ),
    .C1(\adder/adder/_0346_ ),
    .C2(\adder/adder/_0318_ ),
    .ZN(\adder/adder/_0347_ ));
 INV_X1 \adder/adder/_1148_  (.A(\operand_fp16_fp32[24] ),
    .ZN(\adder/adder/_0348_ ));
 NOR2_X1 \adder/adder/_1149_  (.A1(\adder/adder/_0348_ ),
    .A2(net33),
    .ZN(\adder/adder/_0349_ ));
 INV_X1 \adder/adder/_1150_  (.A(\adder/adder/_0349_ ),
    .ZN(\adder/adder/_0350_ ));
 INV_X2 \adder/adder/_1151_  (.A(net33),
    .ZN(\adder/adder/_0351_ ));
 NOR2_X1 \adder/adder/_1152_  (.A1(\adder/adder/_0351_ ),
    .A2(\operand_fp16_fp32[24] ),
    .ZN(\adder/adder/_0352_ ));
 INV_X1 \adder/adder/_1153_  (.A(net32),
    .ZN(\adder/adder/_0353_ ));
 NOR2_X2 \adder/adder/_1154_  (.A1(\adder/adder/_0353_ ),
    .A2(\operand_fp16_fp32[23] ),
    .ZN(\adder/adder/_0354_ ));
 OAI21_X2 \adder/adder/_1155_  (.A(\adder/adder/_0350_ ),
    .B1(\adder/adder/_0352_ ),
    .B2(\adder/adder/_0354_ ),
    .ZN(\adder/adder/_0355_ ));
 INV_X1 \adder/adder/_1156_  (.A(\operand_fp16_fp32[25] ),
    .ZN(\adder/adder/_0356_ ));
 NAND2_X1 \adder/adder/_1157_  (.A1(\adder/adder/_0356_ ),
    .A2(net34),
    .ZN(\adder/adder/_0357_ ));
 INV_X1 \adder/adder/_1158_  (.A(net34),
    .ZN(\adder/adder/_0358_ ));
 NAND2_X1 \adder/adder/_1159_  (.A1(\adder/adder/_0358_ ),
    .A2(\operand_fp16_fp32[25] ),
    .ZN(\adder/adder/_0359_ ));
 NAND2_X1 \adder/adder/_1160_  (.A1(\adder/adder/_0357_ ),
    .A2(\adder/adder/_0359_ ),
    .ZN(\adder/adder/_0360_ ));
 INV_X1 \adder/adder/_1161_  (.A(\adder/adder/_0360_ ),
    .ZN(\adder/adder/_0361_ ));
 NAND2_X1 \adder/adder/_1162_  (.A1(\adder/adder/_0355_ ),
    .A2(\adder/adder/_0361_ ),
    .ZN(\adder/adder/_0362_ ));
 NAND2_X1 \adder/adder/_1163_  (.A1(\adder/adder/_0362_ ),
    .A2(\adder/adder/_0359_ ),
    .ZN(\adder/adder/_0363_ ));
 INV_X1 \adder/adder/_1164_  (.A(\operand_fp16_fp32[26] ),
    .ZN(\adder/adder/_0364_ ));
 NAND2_X1 \adder/adder/_1165_  (.A1(\adder/adder/_0364_ ),
    .A2(net35),
    .ZN(\adder/adder/_0365_ ));
 INV_X1 \adder/adder/_1166_  (.A(net35),
    .ZN(\adder/adder/_0366_ ));
 NAND2_X1 \adder/adder/_1167_  (.A1(\adder/adder/_0366_ ),
    .A2(\operand_fp16_fp32[26] ),
    .ZN(\adder/adder/_0367_ ));
 NAND2_X2 \adder/adder/_1168_  (.A1(\adder/adder/_0365_ ),
    .A2(\adder/adder/_0367_ ),
    .ZN(\adder/adder/_0368_ ));
 INV_X1 \adder/adder/_1169_  (.A(\adder/adder/_0368_ ),
    .ZN(\adder/adder/_0369_ ));
 XNOR2_X1 \adder/adder/_1170_  (.A(\adder/adder/_0363_ ),
    .B(\adder/adder/_0369_ ),
    .ZN(\adder/adder/_0370_ ));
 INV_X1 \adder/adder/_1171_  (.A(\adder/adder/_0352_ ),
    .ZN(\adder/adder/_0371_ ));
 INV_X1 \adder/adder/_1172_  (.A(\operand_fp16_fp32[23] ),
    .ZN(\adder/adder/_0372_ ));
 NOR2_X2 \adder/adder/_1173_  (.A1(\adder/adder/_0372_ ),
    .A2(net32),
    .ZN(\adder/adder/_0373_ ));
 OAI21_X1 \adder/adder/_1174_  (.A(\adder/adder/_0371_ ),
    .B1(\adder/adder/_0373_ ),
    .B2(\adder/adder/_0349_ ),
    .ZN(\adder/adder/_0374_ ));
 NOR2_X2 \adder/adder/_1175_  (.A1(\adder/adder/_0368_ ),
    .A2(\adder/adder/_0360_ ),
    .ZN(\adder/adder/_0375_ ));
 NAND2_X1 \adder/adder/_1176_  (.A1(\adder/adder/_0374_ ),
    .A2(\adder/adder/_0375_ ),
    .ZN(\adder/adder/_0376_ ));
 NOR2_X1 \adder/adder/_1177_  (.A1(\adder/adder/_0368_ ),
    .A2(\adder/adder/_0357_ ),
    .ZN(\adder/adder/_0377_ ));
 INV_X1 \adder/adder/_1178_  (.A(\adder/adder/_0365_ ),
    .ZN(\adder/adder/_0378_ ));
 NOR2_X1 \adder/adder/_1179_  (.A1(\adder/adder/_0377_ ),
    .A2(\adder/adder/_0378_ ),
    .ZN(\adder/adder/_0379_ ));
 NAND2_X2 \adder/adder/_1180_  (.A1(\adder/adder/_0376_ ),
    .A2(\adder/adder/_0379_ ),
    .ZN(\adder/adder/_0380_ ));
 INV_X1 \adder/adder/_1181_  (.A(net6),
    .ZN(\adder/adder/_0381_ ));
 INV_X1 \adder/adder/_1182_  (.A(net40),
    .ZN(\adder/adder/_0382_ ));
 NAND2_X2 \adder/adder/_1183_  (.A1(\adder/adder/_0381_ ),
    .A2(\adder/adder/_0382_ ),
    .ZN(\adder/exp_prenorm_d[7] ));
 NAND2_X1 \adder/adder/_1184_  (.A1(net6),
    .A2(net40),
    .ZN(\adder/adder/_0383_ ));
 NAND2_X1 \adder/adder/_1185_  (.A1(\adder/exp_prenorm_d[7] ),
    .A2(\adder/adder/_0383_ ),
    .ZN(\adder/adder/_0384_ ));
 INV_X2 \adder/adder/_1186_  (.A(\adder/adder/_0384_ ),
    .ZN(\adder/adder/_0385_ ));
 INV_X1 \adder/adder/_1187_  (.A(\operand_fp16_fp32[29] ),
    .ZN(\adder/adder/_0386_ ));
 NAND2_X1 \adder/adder/_1188_  (.A1(\adder/adder/_0386_ ),
    .A2(net38),
    .ZN(\adder/adder/_0387_ ));
 INV_X1 \adder/adder/_1189_  (.A(net38),
    .ZN(\adder/adder/_0388_ ));
 NAND2_X1 \adder/adder/_1190_  (.A1(\adder/adder/_0388_ ),
    .A2(\operand_fp16_fp32[29] ),
    .ZN(\adder/adder/_0389_ ));
 NAND2_X2 \adder/adder/_1191_  (.A1(\adder/adder/_0387_ ),
    .A2(\adder/adder/_0389_ ),
    .ZN(\adder/adder/_0390_ ));
 NOR2_X1 \adder/adder/_1192_  (.A1(\adder/adder/_0385_ ),
    .A2(\adder/adder/_0390_ ),
    .ZN(\adder/adder/_0391_ ));
 INV_X1 \adder/adder/_1193_  (.A(\adder/adder/_0391_ ),
    .ZN(\adder/adder/_0392_ ));
 INV_X2 \adder/adder/_1194_  (.A(\operand_fp16_fp32[27] ),
    .ZN(\adder/adder/_0393_ ));
 NAND2_X1 \adder/adder/_1195_  (.A1(\adder/adder/_0393_ ),
    .A2(net36),
    .ZN(\adder/adder/_0394_ ));
 INV_X1 \adder/adder/_1196_  (.A(\adder/adder/_0394_ ),
    .ZN(\adder/adder/_0395_ ));
 NOR2_X1 \adder/adder/_1197_  (.A1(\adder/adder/_0393_ ),
    .A2(net36),
    .ZN(\adder/adder/_0396_ ));
 NOR2_X2 \adder/adder/_1198_  (.A1(\adder/adder/_0395_ ),
    .A2(\adder/adder/_0396_ ),
    .ZN(\adder/adder/_0397_ ));
 INV_X1 \adder/adder/_1199_  (.A(\operand_fp16_fp32[29] ),
    .ZN(\adder/adder/_0398_ ));
 NAND2_X1 \adder/adder/_1200_  (.A1(\adder/adder/_0398_ ),
    .A2(net37),
    .ZN(\adder/adder/_0399_ ));
 INV_X1 \adder/adder/_1201_  (.A(\adder/adder/_0399_ ),
    .ZN(\adder/adder/_0400_ ));
 NOR2_X1 \adder/adder/_1202_  (.A1(\adder/adder/_0398_ ),
    .A2(net37),
    .ZN(\adder/adder/_0401_ ));
 NOR2_X1 \adder/adder/_1203_  (.A1(\adder/adder/_0400_ ),
    .A2(\adder/adder/_0401_ ),
    .ZN(\adder/adder/_0402_ ));
 NAND2_X1 \adder/adder/_1204_  (.A1(\adder/adder/_0397_ ),
    .A2(\adder/adder/_0402_ ),
    .ZN(\adder/adder/_0403_ ));
 NOR2_X1 \adder/adder/_1205_  (.A1(\adder/adder/_0392_ ),
    .A2(\adder/adder/_0403_ ),
    .ZN(\adder/adder/_0404_ ));
 NAND2_X2 \adder/adder/_1206_  (.A1(\adder/adder/_0380_ ),
    .A2(\adder/adder/_0404_ ),
    .ZN(\adder/adder/_0405_ ));
 OAI21_X1 \adder/adder/_1207_  (.A(\adder/adder/_0399_ ),
    .B1(\adder/adder/_0401_ ),
    .B2(\adder/adder/_0394_ ),
    .ZN(\adder/adder/_0406_ ));
 NAND2_X1 \adder/adder/_1208_  (.A1(\adder/adder/_0391_ ),
    .A2(\adder/adder/_0406_ ),
    .ZN(\adder/adder/_0407_ ));
 NOR2_X1 \adder/adder/_1209_  (.A1(\adder/adder/_0382_ ),
    .A2(net6),
    .ZN(\adder/adder/_0408_ ));
 INV_X1 \adder/adder/_1210_  (.A(\adder/adder/_0387_ ),
    .ZN(\adder/adder/_0409_ ));
 AOI21_X1 \adder/adder/_1211_  (.A(\adder/adder/_0408_ ),
    .B1(\adder/adder/_0384_ ),
    .B2(\adder/adder/_0409_ ),
    .ZN(\adder/adder/_0410_ ));
 NAND2_X1 \adder/adder/_1212_  (.A1(\adder/adder/_0407_ ),
    .A2(\adder/adder/_0410_ ),
    .ZN(\adder/adder/_0411_ ));
 INV_X1 \adder/adder/_1213_  (.A(\adder/adder/_0411_ ),
    .ZN(\adder/adder/_0412_ ));
 NAND2_X4 \adder/adder/_1214_  (.A1(\adder/adder/_0412_ ),
    .A2(\adder/adder/_0405_ ),
    .ZN(\adder/adder/_0413_ ));
 INV_X8 \adder/adder/_1215_  (.A(\adder/adder/_0413_ ),
    .ZN(\adder/adder/_0414_ ));
 NAND2_X1 \adder/adder/_1216_  (.A1(\adder/adder/_0370_ ),
    .A2(\adder/adder/_0414_ ),
    .ZN(\adder/adder/_0415_ ));
 NAND2_X1 \adder/adder/_1217_  (.A1(\adder/adder/_0374_ ),
    .A2(\adder/adder/_0361_ ),
    .ZN(\adder/adder/_0416_ ));
 NAND2_X1 \adder/adder/_1218_  (.A1(\adder/adder/_0416_ ),
    .A2(\adder/adder/_0357_ ),
    .ZN(\adder/adder/_0417_ ));
 XNOR2_X1 \adder/adder/_1219_  (.A(\adder/adder/_0417_ ),
    .B(\adder/adder/_0369_ ),
    .ZN(\adder/adder/_0418_ ));
 NAND2_X1 \adder/adder/_1220_  (.A1(\adder/adder/_0418_ ),
    .A2(\adder/adder/_0413_ ),
    .ZN(\adder/adder/_0419_ ));
 NAND2_X4 \adder/adder/_1221_  (.A1(\adder/adder/_0419_ ),
    .A2(\adder/adder/_0415_ ),
    .ZN(\adder/adder/_0420_ ));
 INV_X16 \adder/adder/_1222_  (.A(\adder/adder/_0420_ ),
    .ZN(\adder/adder/_0421_ ));
 BUF_X16 max_cap83 (.A(net84),
    .Z(net83));
 NOR2_X1 \adder/adder/_1224_  (.A1(\adder/adder/_0347_ ),
    .A2(\adder/adder/_0421_ ),
    .ZN(\adder/adder/_0423_ ));
 NAND2_X1 \adder/adder/_1225_  (.A1(\adder/adder/_0355_ ),
    .A2(\adder/adder/_0375_ ),
    .ZN(\adder/adder/_0424_ ));
 NOR2_X1 \adder/adder/_1226_  (.A1(\adder/adder/_0368_ ),
    .A2(\adder/adder/_0359_ ),
    .ZN(\adder/adder/_0425_ ));
 INV_X1 \adder/adder/_1227_  (.A(\adder/adder/_0367_ ),
    .ZN(\adder/adder/_0426_ ));
 NOR2_X1 \adder/adder/_1228_  (.A1(\adder/adder/_0425_ ),
    .A2(\adder/adder/_0426_ ),
    .ZN(\adder/adder/_0427_ ));
 NAND2_X1 \adder/adder/_1229_  (.A1(\adder/adder/_0424_ ),
    .A2(\adder/adder/_0427_ ),
    .ZN(\adder/adder/_0428_ ));
 AOI21_X1 \adder/adder/_1230_  (.A(\adder/adder/_0396_ ),
    .B1(\adder/adder/_0428_ ),
    .B2(\adder/adder/_0397_ ),
    .ZN(\adder/adder/_0429_ ));
 NAND2_X1 \adder/adder/_1231_  (.A1(\adder/adder/_0414_ ),
    .A2(\adder/adder/_0429_ ),
    .ZN(\adder/adder/_0430_ ));
 AOI21_X1 \adder/adder/_1232_  (.A(\adder/adder/_0395_ ),
    .B1(\adder/adder/_0380_ ),
    .B2(\adder/adder/_0397_ ),
    .ZN(\adder/adder/_0431_ ));
 NAND2_X1 \adder/adder/_1233_  (.A1(\adder/adder/_0431_ ),
    .A2(\adder/adder/_0413_ ),
    .ZN(\adder/adder/_0432_ ));
 NAND2_X1 \adder/adder/_1234_  (.A1(\adder/adder/_0430_ ),
    .A2(\adder/adder/_0432_ ),
    .ZN(\adder/adder/_0433_ ));
 OAI21_X1 \adder/adder/_1235_  (.A(\adder/adder/_0433_ ),
    .B1(\adder/adder/_0400_ ),
    .B2(\adder/adder/_0401_ ),
    .ZN(\adder/adder/_0434_ ));
 NAND3_X1 \adder/adder/_1236_  (.A1(\adder/adder/_0430_ ),
    .A2(\adder/adder/_0432_ ),
    .A3(\adder/adder/_0402_ ),
    .ZN(\adder/adder/_0435_ ));
 NAND2_X2 \adder/adder/_1237_  (.A1(\adder/adder/_0434_ ),
    .A2(\adder/adder/_0435_ ),
    .ZN(\adder/adder/_0436_ ));
 INV_X2 \adder/adder/_1238_  (.A(\adder/adder/_0436_ ),
    .ZN(\adder/adder/_0437_ ));
 XOR2_X1 \adder/adder/_1239_  (.A(\adder/adder/_0380_ ),
    .B(\adder/adder/_0397_ ),
    .Z(\adder/adder/_0438_ ));
 NAND2_X1 \adder/adder/_1240_  (.A1(\adder/adder/_0438_ ),
    .A2(\adder/adder/_0413_ ),
    .ZN(\adder/adder/_0439_ ));
 XOR2_X1 \adder/adder/_1241_  (.A(\adder/adder/_0428_ ),
    .B(\adder/adder/_0397_ ),
    .Z(\adder/adder/_0440_ ));
 NAND2_X1 \adder/adder/_1242_  (.A1(\adder/adder/_0440_ ),
    .A2(\adder/adder/_0414_ ),
    .ZN(\adder/adder/_0441_ ));
 NAND2_X2 \adder/adder/_1243_  (.A1(\adder/adder/_0439_ ),
    .A2(\adder/adder/_0441_ ),
    .ZN(\adder/adder/_0442_ ));
 NOR2_X4 \adder/adder/_1244_  (.A1(\adder/adder/_0442_ ),
    .A2(\adder/adder/_0437_ ),
    .ZN(\adder/adder/_0443_ ));
 NAND2_X1 \adder/adder/_1245_  (.A1(\adder/adder/_0371_ ),
    .A2(\adder/adder/_0350_ ),
    .ZN(\adder/adder/_0444_ ));
 XNOR2_X1 \adder/adder/_1246_  (.A(\adder/adder/_0444_ ),
    .B(\adder/adder/_0373_ ),
    .ZN(\adder/adder/_0445_ ));
 NAND2_X1 \adder/adder/_1247_  (.A1(\adder/adder/_0413_ ),
    .A2(\adder/adder/_0445_ ),
    .ZN(\adder/adder/_0446_ ));
 XNOR2_X1 \adder/adder/_1248_  (.A(\adder/adder/_0444_ ),
    .B(\adder/adder/_0354_ ),
    .ZN(\adder/adder/_0447_ ));
 NAND3_X2 \adder/adder/_1249_  (.A1(\adder/adder/_0405_ ),
    .A2(\adder/adder/_0412_ ),
    .A3(\adder/adder/_0447_ ),
    .ZN(\adder/adder/_0448_ ));
 NAND2_X4 \adder/adder/_1250_  (.A1(\adder/adder/_0448_ ),
    .A2(\adder/adder/_0446_ ),
    .ZN(\adder/adder/_0449_ ));
 INV_X4 \adder/adder/_1251_  (.A(\adder/adder/_0449_ ),
    .ZN(\adder/adder/_0450_ ));
 NOR2_X4 \adder/adder/_1252_  (.A1(\adder/adder/_0373_ ),
    .A2(\adder/adder/_0354_ ),
    .ZN(\adder/adder/_0451_ ));
 INV_X8 \adder/adder/_1253_  (.A(\adder/adder/_0451_ ),
    .ZN(\adder/adder/_0452_ ));
 NOR2_X1 \adder/adder/_1254_  (.A1(\adder/adder/_0450_ ),
    .A2(\adder/adder/_0452_ ),
    .ZN(\adder/adder/_0453_ ));
 XNOR2_X1 \adder/adder/_1255_  (.A(\adder/adder/_0355_ ),
    .B(\adder/adder/_0361_ ),
    .ZN(\adder/adder/_0454_ ));
 NAND2_X1 \adder/adder/_1256_  (.A1(\adder/adder/_0414_ ),
    .A2(\adder/adder/_0454_ ),
    .ZN(\adder/adder/_0455_ ));
 XNOR2_X1 \adder/adder/_1257_  (.A(\adder/adder/_0374_ ),
    .B(\adder/adder/_0361_ ),
    .ZN(\adder/adder/_0456_ ));
 NAND2_X1 \adder/adder/_1258_  (.A1(\adder/adder/_0413_ ),
    .A2(\adder/adder/_0456_ ),
    .ZN(\adder/adder/_0457_ ));
 NAND2_X4 \adder/adder/_1259_  (.A1(\adder/adder/_0457_ ),
    .A2(\adder/adder/_0455_ ),
    .ZN(\adder/adder/_0458_ ));
 NAND4_X1 \adder/adder/_1260_  (.A1(\adder/adder/_0423_ ),
    .A2(\adder/adder/_0443_ ),
    .A3(\adder/adder/_0453_ ),
    .A4(\adder/adder/_0458_ ),
    .ZN(\adder/adder/_0459_ ));
 INV_X1 \adder/adder/_1261_  (.A(\adder/adder/_0403_ ),
    .ZN(\adder/adder/_0460_ ));
 AOI21_X1 \adder/adder/_1262_  (.A(\adder/adder/_0406_ ),
    .B1(\adder/adder/_0380_ ),
    .B2(\adder/adder/_0460_ ),
    .ZN(\adder/adder/_0461_ ));
 NAND2_X1 \adder/adder/_1263_  (.A1(\adder/adder/_0461_ ),
    .A2(\adder/adder/_0413_ ),
    .ZN(\adder/adder/_0462_ ));
 NAND2_X1 \adder/adder/_1264_  (.A1(\adder/adder/_0428_ ),
    .A2(\adder/adder/_0460_ ),
    .ZN(\adder/adder/_0463_ ));
 AOI21_X1 \adder/adder/_1265_  (.A(\adder/adder/_0401_ ),
    .B1(\adder/adder/_0399_ ),
    .B2(\adder/adder/_0396_ ),
    .ZN(\adder/adder/_0464_ ));
 NAND2_X1 \adder/adder/_1266_  (.A1(\adder/adder/_0463_ ),
    .A2(\adder/adder/_0464_ ),
    .ZN(\adder/adder/_0465_ ));
 OAI21_X1 \adder/adder/_1267_  (.A(\adder/adder/_0462_ ),
    .B1(\adder/adder/_0413_ ),
    .B2(\adder/adder/_0465_ ),
    .ZN(\adder/adder/_0466_ ));
 XNOR2_X2 \adder/adder/_1268_  (.A(\adder/adder/_0466_ ),
    .B(\adder/adder/_0390_ ),
    .ZN(\adder/adder/_0467_ ));
 NOR2_X1 \adder/adder/_1269_  (.A1(\adder/adder/_0414_ ),
    .A2(\adder/adder/_0409_ ),
    .ZN(\adder/adder/_0468_ ));
 OAI21_X1 \adder/adder/_1270_  (.A(\adder/adder/_0468_ ),
    .B1(\adder/adder/_0390_ ),
    .B2(\adder/adder/_0461_ ),
    .ZN(\adder/adder/_0469_ ));
 INV_X1 \adder/adder/_1271_  (.A(\adder/adder/_0390_ ),
    .ZN(\adder/adder/_0470_ ));
 NAND2_X1 \adder/adder/_1272_  (.A1(\adder/adder/_0465_ ),
    .A2(\adder/adder/_0470_ ),
    .ZN(\adder/adder/_0471_ ));
 NAND3_X2 \adder/adder/_1273_  (.A1(\adder/adder/_0471_ ),
    .A2(\adder/adder/_0389_ ),
    .A3(\adder/adder/_0414_ ),
    .ZN(\adder/adder/_0472_ ));
 NAND3_X4 \adder/adder/_1274_  (.A1(\adder/adder/_0469_ ),
    .A2(\adder/adder/_0385_ ),
    .A3(\adder/adder/_0472_ ),
    .ZN(\adder/adder/_0473_ ));
 NAND2_X4 \adder/adder/_1275_  (.A1(\adder/adder/_0467_ ),
    .A2(\adder/adder/_0473_ ),
    .ZN(\adder/adder/_0474_ ));
 BUF_X16 max_cap82 (.A(\adder/norm/_0680_ ),
    .Z(net82));
 NOR2_X2 \adder/adder/_1277_  (.A1(\adder/adder/_0459_ ),
    .A2(\adder/adder/_0474_ ),
    .ZN(\adder/adder/_0476_ ));
 NAND2_X2 \adder/adder/_1278_  (.A1(\adder/adder/_0337_ ),
    .A2(\adder/adder/_0476_ ),
    .ZN(\adder/adder/_0477_ ));
 BUF_X16 max_cap81 (.A(net82),
    .Z(net81));
 BUF_X1 output80 (.A(net80),
    .Z(result_o[9]));
 BUF_X1 output79 (.A(net79),
    .Z(result_o[8]));
 BUF_X1 output78 (.A(net78),
    .Z(result_o[7]));
 BUF_X1 output77 (.A(net77),
    .Z(result_o[6]));
 BUF_X1 output76 (.A(net76),
    .Z(result_o[5]));
 BUF_X1 output75 (.A(net75),
    .Z(result_o[4]));
 NAND2_X1 \adder/adder/_1286_  (.A1(\adder/adder/_0477_ ),
    .A2(net239),
    .ZN(\adder/adder/_0485_ ));
 MUX2_X1 \adder/adder/_1287_  (.A(net41),
    .B(net7),
    .S(\adder/adder/_0485_ ),
    .Z(net73));
 BUF_X1 output74 (.A(net74),
    .Z(result_o[3]));
 NAND2_X1 \adder/adder/_1289_  (.A1(net239),
    .A2(net32),
    .ZN(\adder/adder/_0487_ ));
 OAI21_X2 \adder/adder/_1290_  (.A(\adder/adder/_0487_ ),
    .B1(\adder/adder/_0372_ ),
    .B2(net239),
    .ZN(\adder/exp_prenorm_d[0] ));
 NAND2_X1 \adder/adder/_1291_  (.A1(net239),
    .A2(net33),
    .ZN(\adder/adder/_0488_ ));
 OAI21_X1 \adder/adder/_1292_  (.A(\adder/adder/_0488_ ),
    .B1(\adder/adder/_0348_ ),
    .B2(net239),
    .ZN(\adder/exp_prenorm_d[1] ));
 NAND2_X1 \adder/adder/_1293_  (.A1(net239),
    .A2(net34),
    .ZN(\adder/adder/_0489_ ));
 OAI21_X1 \adder/adder/_1294_  (.A(\adder/adder/_0489_ ),
    .B1(\adder/adder/_0356_ ),
    .B2(net239),
    .ZN(\adder/exp_prenorm_d[2] ));
 NAND2_X1 \adder/adder/_1295_  (.A1(net239),
    .A2(net35),
    .ZN(\adder/adder/_0490_ ));
 OAI21_X1 \adder/adder/_1296_  (.A(\adder/adder/_0490_ ),
    .B1(\adder/adder/_0364_ ),
    .B2(net239),
    .ZN(\adder/exp_prenorm_d[3] ));
 NAND2_X1 \adder/adder/_1297_  (.A1(net239),
    .A2(net36),
    .ZN(\adder/adder/_0491_ ));
 OAI21_X1 \adder/adder/_1298_  (.A(\adder/adder/_0491_ ),
    .B1(\adder/adder/_0393_ ),
    .B2(net239),
    .ZN(\adder/exp_prenorm_d[4] ));
 NAND2_X1 \adder/adder/_1299_  (.A1(net239),
    .A2(net37),
    .ZN(\adder/adder/_0492_ ));
 OAI21_X2 \adder/adder/_1300_  (.A(\adder/adder/_0492_ ),
    .B1(\adder/adder/_0398_ ),
    .B2(net239),
    .ZN(\adder/exp_prenorm_d[5] ));
 NAND2_X1 \adder/adder/_1301_  (.A1(net239),
    .A2(net38),
    .ZN(\adder/adder/_0493_ ));
 OAI21_X2 \adder/adder/_1302_  (.A(\adder/adder/_0493_ ),
    .B1(\adder/adder/_0386_ ),
    .B2(net239),
    .ZN(\adder/exp_prenorm_d[6] ));
 XNOR2_X2 \adder/adder/_1303_  (.A(net7),
    .B(net41),
    .ZN(\adder/adder/_0494_ ));
 INV_X2 \adder/adder/_1304_  (.A(\adder/adder/_0494_ ),
    .ZN(\adder/adder/_0495_ ));
 NAND3_X1 \adder/adder/_1305_  (.A1(\adder/adder/_0446_ ),
    .A2(\adder/adder/_0448_ ),
    .A3(\adder/adder/_0452_ ),
    .ZN(\adder/adder/_0496_ ));
 INV_X1 \adder/adder/_1306_  (.A(\adder/adder/_0496_ ),
    .ZN(\adder/adder/_0497_ ));
 INV_X4 \adder/adder/_1307_  (.A(\adder/adder/_0458_ ),
    .ZN(\adder/adder/_0498_ ));
 NAND2_X1 \adder/adder/_1308_  (.A1(\adder/adder/_0497_ ),
    .A2(\adder/adder/_0498_ ),
    .ZN(\adder/adder/_0499_ ));
 NAND2_X2 \adder/adder/_1309_  (.A1(\adder/adder/_0496_ ),
    .A2(\adder/adder/_0458_ ),
    .ZN(\adder/adder/_0500_ ));
 AND2_X1 \adder/adder/_1310_  (.A1(\adder/adder/_0499_ ),
    .A2(\adder/adder/_0500_ ),
    .ZN(\adder/adder/_0501_ ));
 NAND3_X2 \adder/adder/_1311_  (.A1(\adder/adder/_0500_ ),
    .A2(\adder/adder/_0442_ ),
    .A3(\adder/adder/_0421_ ),
    .ZN(\adder/adder/_0502_ ));
 NAND2_X2 \adder/adder/_1312_  (.A1(\adder/adder/_0502_ ),
    .A2(\adder/adder/_0436_ ),
    .ZN(\adder/adder/_0503_ ));
 INV_X1 \adder/adder/_1313_  (.A(\adder/adder/_0467_ ),
    .ZN(\adder/adder/_0504_ ));
 NAND2_X1 \adder/adder/_1314_  (.A1(\adder/adder/_0503_ ),
    .A2(\adder/adder/_0504_ ),
    .ZN(\adder/adder/_0505_ ));
 NAND2_X4 \adder/adder/_1315_  (.A1(\adder/adder/_0474_ ),
    .A2(\adder/adder/_0505_ ),
    .ZN(\adder/adder/_0506_ ));
 BUF_X1 output73 (.A(net73),
    .Z(result_o[31]));
 NAND2_X1 \adder/adder/_1317_  (.A1(net239),
    .A2(net202),
    .ZN(\adder/adder/_0508_ ));
 BUF_X1 output72 (.A(net72),
    .Z(result_o[30]));
 OAI21_X1 \adder/adder/_1319_  (.A(\adder/adder/_0508_ ),
    .B1(\adder/adder/_0266_ ),
    .B2(net242),
    .ZN(\adder/adder/_0510_ ));
 NAND2_X4 \adder/adder/_1320_  (.A1(\adder/adder/_0503_ ),
    .A2(\adder/adder/_0473_ ),
    .ZN(\adder/adder/_0511_ ));
 BUF_X1 output71 (.A(net71),
    .Z(result_o[2]));
 NAND3_X1 \adder/adder/_1322_  (.A1(\adder/adder/_0506_ ),
    .A2(\adder/adder/_0510_ ),
    .A3(\adder/adder/_0511_ ),
    .ZN(\adder/adder/_0513_ ));
 BUF_X1 output70 (.A(net70),
    .Z(result_o[29]));
 BUF_X1 output69 (.A(net69),
    .Z(result_o[28]));
 NAND2_X1 \adder/adder/_1325_  (.A1(\adder/adder/_0513_ ),
    .A2(\adder/adder/_0452_ ),
    .ZN(\adder/adder/_0516_ ));
 NAND2_X1 \adder/adder/_1326_  (.A1(net242),
    .A2(\adder/adder/_0261_ ),
    .ZN(\adder/adder/_0517_ ));
 BUF_X1 output68 (.A(net68),
    .Z(result_o[27]));
 OAI21_X1 \adder/adder/_1328_  (.A(\adder/adder/_0517_ ),
    .B1(net20),
    .B2(net245),
    .ZN(\adder/adder/_0519_ ));
 INV_X1 \adder/adder/_1329_  (.A(\adder/adder/_0519_ ),
    .ZN(\adder/adder/_0520_ ));
 NAND3_X1 \adder/adder/_1330_  (.A1(\adder/adder/_0506_ ),
    .A2(\adder/adder/_0520_ ),
    .A3(\adder/adder/_0511_ ),
    .ZN(\adder/adder/_0521_ ));
 BUF_X1 output67 (.A(net67),
    .Z(result_o[26]));
 BUF_X1 output66 (.A(net66),
    .Z(result_o[25]));
 NAND2_X1 \adder/adder/_1333_  (.A1(\adder/adder/_0521_ ),
    .A2(\adder/adder/_0451_ ),
    .ZN(\adder/adder/_0524_ ));
 NAND2_X1 \adder/adder/_1334_  (.A1(\adder/adder/_0516_ ),
    .A2(\adder/adder/_0524_ ),
    .ZN(\adder/adder/_0525_ ));
 BUF_X1 output65 (.A(net65),
    .Z(result_o[24]));
 NAND2_X1 \adder/adder/_1336_  (.A1(\adder/adder/_0521_ ),
    .A2(\adder/adder/_0452_ ),
    .ZN(\adder/adder/_0527_ ));
 BUF_X1 output64 (.A(net64),
    .Z(result_o[23]));
 NAND2_X1 \adder/adder/_1338_  (.A1(\adder/adder/_0414_ ),
    .A2(\adder/adder/_0284_ ),
    .ZN(\adder/adder/_0529_ ));
 OAI21_X1 \adder/adder/_1339_  (.A(\adder/adder/_0529_ ),
    .B1(\operand_fp16_fp32[13] ),
    .B2(\adder/adder/_0414_ ),
    .ZN(\adder/adder/_0530_ ));
 INV_X1 \adder/adder/_1340_  (.A(\adder/adder/_0530_ ),
    .ZN(\adder/adder/_0531_ ));
 NAND3_X1 \adder/adder/_1341_  (.A1(\adder/adder/_0506_ ),
    .A2(\adder/adder/_0531_ ),
    .A3(\adder/adder/_0511_ ),
    .ZN(\adder/adder/_0532_ ));
 BUF_X1 output63 (.A(net63),
    .Z(result_o[22]));
 BUF_X1 output62 (.A(net62),
    .Z(result_o[21]));
 NAND2_X1 \adder/adder/_1344_  (.A1(\adder/adder/_0532_ ),
    .A2(\adder/adder/_0451_ ),
    .ZN(\adder/adder/_0535_ ));
 NAND2_X1 \adder/adder/_1345_  (.A1(\adder/adder/_0527_ ),
    .A2(\adder/adder/_0535_ ),
    .ZN(\adder/adder/_0536_ ));
 OR2_X4 \adder/adder/_1346_  (.A1(\adder/adder/_0453_ ),
    .A2(\adder/adder/_0497_ ),
    .ZN(\adder/adder/_0537_ ));
 INV_X2 \adder/adder/_1347_  (.A(\adder/adder/_0537_ ),
    .ZN(\adder/adder/_0538_ ));
 NAND3_X1 \adder/adder/_1348_  (.A1(\adder/adder/_0525_ ),
    .A2(\adder/adder/_0536_ ),
    .A3(\adder/adder/_0538_ ),
    .ZN(\adder/adder/_0539_ ));
 NAND2_X1 \adder/adder/_1349_  (.A1(net245),
    .A2(\adder/adder/_0270_ ),
    .ZN(\adder/adder/_0540_ ));
 OAI21_X1 \adder/adder/_1350_  (.A(\adder/adder/_0540_ ),
    .B1(net18),
    .B2(net245),
    .ZN(\adder/adder/_0541_ ));
 INV_X1 \adder/adder/_1351_  (.A(\adder/adder/_0541_ ),
    .ZN(\adder/adder/_0542_ ));
 NAND3_X1 \adder/adder/_1352_  (.A1(\adder/adder/_0506_ ),
    .A2(\adder/adder/_0542_ ),
    .A3(\adder/adder/_0511_ ),
    .ZN(\adder/adder/_0543_ ));
 NAND2_X1 \adder/adder/_1353_  (.A1(\adder/adder/_0543_ ),
    .A2(\adder/adder/_0452_ ),
    .ZN(\adder/adder/_0544_ ));
 NAND2_X1 \adder/adder/_1354_  (.A1(\adder/adder/_0513_ ),
    .A2(\adder/adder/_0451_ ),
    .ZN(\adder/adder/_0545_ ));
 NAND2_X1 \adder/adder/_1355_  (.A1(\adder/adder/_0544_ ),
    .A2(\adder/adder/_0545_ ),
    .ZN(\adder/adder/_0546_ ));
 OR2_X1 \adder/adder/_1356_  (.A1(\adder/adder/_0414_ ),
    .A2(net203),
    .ZN(\adder/adder/_0547_ ));
 OAI21_X1 \adder/adder/_1357_  (.A(\adder/adder/_0547_ ),
    .B1(net48),
    .B2(net245),
    .ZN(\adder/adder/_0548_ ));
 INV_X1 \adder/adder/_1358_  (.A(\adder/adder/_0548_ ),
    .ZN(\adder/adder/_0549_ ));
 NAND3_X1 \adder/adder/_1359_  (.A1(\adder/adder/_0506_ ),
    .A2(\adder/adder/_0549_ ),
    .A3(\adder/adder/_0511_ ),
    .ZN(\adder/adder/_0550_ ));
 NAND2_X1 \adder/adder/_1360_  (.A1(\adder/adder/_0550_ ),
    .A2(\adder/adder/_0452_ ),
    .ZN(\adder/adder/_0551_ ));
 NAND2_X1 \adder/adder/_1361_  (.A1(\adder/adder/_0543_ ),
    .A2(net85),
    .ZN(\adder/adder/_0552_ ));
 NAND2_X1 \adder/adder/_1362_  (.A1(\adder/adder/_0551_ ),
    .A2(\adder/adder/_0552_ ),
    .ZN(\adder/adder/_0553_ ));
 BUF_X1 output61 (.A(net61),
    .Z(result_o[20]));
 NAND3_X1 \adder/adder/_1364_  (.A1(\adder/adder/_0546_ ),
    .A2(\adder/adder/_0553_ ),
    .A3(\adder/adder/_0537_ ),
    .ZN(\adder/adder/_0555_ ));
 NAND2_X1 \adder/adder/_1365_  (.A1(\adder/adder/_0539_ ),
    .A2(\adder/adder/_0555_ ),
    .ZN(\adder/adder/_0556_ ));
 NAND2_X1 \adder/adder/_1366_  (.A1(net242),
    .A2(\operand_fp16_fp32[14] ),
    .ZN(\adder/adder/_0557_ ));
 OAI21_X2 \adder/adder/_1367_  (.A(\adder/adder/_0557_ ),
    .B1(\adder/adder/_0253_ ),
    .B2(net242),
    .ZN(\adder/adder/_0558_ ));
 NAND3_X1 \adder/adder/_1368_  (.A1(\adder/adder/_0506_ ),
    .A2(\adder/adder/_0558_ ),
    .A3(\adder/adder/_0511_ ),
    .ZN(\adder/adder/_0559_ ));
 NAND2_X1 \adder/adder/_1369_  (.A1(\adder/adder/_0559_ ),
    .A2(\adder/adder/_0452_ ),
    .ZN(\adder/adder/_0560_ ));
 BUF_X1 output60 (.A(net60),
    .Z(result_o[1]));
 NAND2_X1 \adder/adder/_1371_  (.A1(net242),
    .A2(\adder/adder/_0255_ ),
    .ZN(\adder/adder/_0562_ ));
 OAI21_X1 \adder/adder/_1372_  (.A(\adder/adder/_0562_ ),
    .B1(net23),
    .B2(net242),
    .ZN(\adder/adder/_0563_ ));
 INV_X1 \adder/adder/_1373_  (.A(\adder/adder/_0563_ ),
    .ZN(\adder/adder/_0564_ ));
 BUF_X1 output59 (.A(net59),
    .Z(result_o[19]));
 NAND3_X1 \adder/adder/_1375_  (.A1(net255),
    .A2(\adder/adder/_0564_ ),
    .A3(\adder/adder/_0511_ ),
    .ZN(\adder/adder/_0566_ ));
 BUF_X1 output58 (.A(net58),
    .Z(result_o[18]));
 NAND2_X1 \adder/adder/_1377_  (.A1(\adder/adder/_0566_ ),
    .A2(\adder/adder/_0451_ ),
    .ZN(\adder/adder/_0568_ ));
 NAND2_X1 \adder/adder/_1378_  (.A1(\adder/adder/_0560_ ),
    .A2(\adder/adder/_0568_ ),
    .ZN(\adder/adder/_0569_ ));
 NAND2_X1 \adder/adder/_1379_  (.A1(\adder/adder/_0532_ ),
    .A2(\adder/adder/_0452_ ),
    .ZN(\adder/adder/_0570_ ));
 NAND2_X1 \adder/adder/_1380_  (.A1(\adder/adder/_0559_ ),
    .A2(\adder/adder/_0451_ ),
    .ZN(\adder/adder/_0571_ ));
 NAND2_X1 \adder/adder/_1381_  (.A1(\adder/adder/_0570_ ),
    .A2(\adder/adder/_0571_ ),
    .ZN(\adder/adder/_0572_ ));
 NAND3_X1 \adder/adder/_1382_  (.A1(\adder/adder/_0569_ ),
    .A2(\adder/adder/_0572_ ),
    .A3(\adder/adder/_0537_ ),
    .ZN(\adder/adder/_0573_ ));
 NAND2_X1 \adder/adder/_1383_  (.A1(net251),
    .A2(\adder/adder/_0333_ ),
    .ZN(\adder/adder/_0574_ ));
 OAI21_X1 \adder/adder/_1384_  (.A(\adder/adder/_0574_ ),
    .B1(net24),
    .B2(net245),
    .ZN(\adder/adder/_0575_ ));
 INV_X1 \adder/adder/_1385_  (.A(\adder/adder/_0575_ ),
    .ZN(\adder/adder/_0576_ ));
 NAND3_X1 \adder/adder/_1386_  (.A1(\adder/adder/_0506_ ),
    .A2(\adder/adder/_0576_ ),
    .A3(\adder/adder/_0511_ ),
    .ZN(\adder/adder/_0577_ ));
 NAND2_X1 \adder/adder/_1387_  (.A1(\adder/adder/_0577_ ),
    .A2(\adder/adder/_0452_ ),
    .ZN(\adder/adder/_0578_ ));
 NAND2_X1 \adder/adder/_1388_  (.A1(net245),
    .A2(\adder/adder/_0319_ ),
    .ZN(\adder/adder/_0579_ ));
 OAI21_X1 \adder/adder/_1389_  (.A(\adder/adder/_0579_ ),
    .B1(net25),
    .B2(net245),
    .ZN(\adder/adder/_0580_ ));
 INV_X1 \adder/adder/_1390_  (.A(\adder/adder/_0580_ ),
    .ZN(\adder/adder/_0581_ ));
 NAND3_X1 \adder/adder/_1391_  (.A1(\adder/adder/_0506_ ),
    .A2(\adder/adder/_0581_ ),
    .A3(\adder/adder/_0511_ ),
    .ZN(\adder/adder/_0582_ ));
 NAND2_X1 \adder/adder/_1392_  (.A1(\adder/adder/_0582_ ),
    .A2(\adder/adder/_0451_ ),
    .ZN(\adder/adder/_0583_ ));
 NAND2_X1 \adder/adder/_1393_  (.A1(\adder/adder/_0578_ ),
    .A2(\adder/adder/_0583_ ),
    .ZN(\adder/adder/_0584_ ));
 NAND2_X1 \adder/adder/_1394_  (.A1(\adder/adder/_0582_ ),
    .A2(\adder/adder/_0452_ ),
    .ZN(\adder/adder/_0585_ ));
 NAND2_X1 \adder/adder/_1395_  (.A1(net242),
    .A2(\operand_fp16_fp32[18] ),
    .ZN(\adder/adder/_0586_ ));
 OAI21_X2 \adder/adder/_1396_  (.A(\adder/adder/_0586_ ),
    .B1(\adder/adder/_0326_ ),
    .B2(net242),
    .ZN(\adder/adder/_0587_ ));
 NAND3_X1 \adder/adder/_1397_  (.A1(\adder/adder/_0506_ ),
    .A2(\adder/adder/_0587_ ),
    .A3(\adder/adder/_0511_ ),
    .ZN(\adder/adder/_0588_ ));
 NAND2_X1 \adder/adder/_1398_  (.A1(\adder/adder/_0588_ ),
    .A2(\adder/adder/_0451_ ),
    .ZN(\adder/adder/_0589_ ));
 NAND2_X1 \adder/adder/_1399_  (.A1(\adder/adder/_0585_ ),
    .A2(\adder/adder/_0589_ ),
    .ZN(\adder/adder/_0590_ ));
 NAND3_X1 \adder/adder/_1400_  (.A1(\adder/adder/_0584_ ),
    .A2(\adder/adder/_0590_ ),
    .A3(\adder/adder/_0538_ ),
    .ZN(\adder/adder/_0591_ ));
 NAND2_X1 \adder/adder/_1401_  (.A1(\adder/adder/_0573_ ),
    .A2(\adder/adder/_0591_ ),
    .ZN(\adder/adder/_0592_ ));
 NAND2_X1 \adder/adder/_1402_  (.A1(\adder/adder/_0556_ ),
    .A2(\adder/adder/_0592_ ),
    .ZN(\adder/adder/_0593_ ));
 NAND2_X1 \adder/adder/_1403_  (.A1(\adder/adder/_0572_ ),
    .A2(\adder/adder/_0538_ ),
    .ZN(\adder/adder/_0594_ ));
 NAND2_X1 \adder/adder/_1404_  (.A1(\adder/adder/_0525_ ),
    .A2(\adder/adder/_0537_ ),
    .ZN(\adder/adder/_0595_ ));
 NAND2_X1 \adder/adder/_1405_  (.A1(\adder/adder/_0594_ ),
    .A2(\adder/adder/_0595_ ),
    .ZN(\adder/adder/_0596_ ));
 NAND4_X1 \adder/adder/_1406_  (.A1(net255),
    .A2(\adder/adder/_0451_ ),
    .A3(\adder/adder/_0564_ ),
    .A4(\adder/adder/_0511_ ),
    .ZN(\adder/adder/_0597_ ));
 NAND4_X1 \adder/adder/_1407_  (.A1(net255),
    .A2(\adder/adder/_0452_ ),
    .A3(\adder/adder/_0558_ ),
    .A4(\adder/adder/_0511_ ),
    .ZN(\adder/adder/_0598_ ));
 NAND3_X1 \adder/adder/_1408_  (.A1(\adder/adder/_0597_ ),
    .A2(\adder/adder/_0598_ ),
    .A3(\adder/adder/_0538_ ),
    .ZN(\adder/adder/_0599_ ));
 NAND4_X1 \adder/adder/_1409_  (.A1(net255),
    .A2(\adder/adder/_0451_ ),
    .A3(\adder/adder/_0531_ ),
    .A4(\adder/adder/_0511_ ),
    .ZN(\adder/adder/_0600_ ));
 NAND4_X1 \adder/adder/_1410_  (.A1(net255),
    .A2(\adder/adder/_0452_ ),
    .A3(\adder/adder/_0520_ ),
    .A4(\adder/adder/_0511_ ),
    .ZN(\adder/adder/_0601_ ));
 NAND3_X1 \adder/adder/_1411_  (.A1(\adder/adder/_0600_ ),
    .A2(\adder/adder/_0601_ ),
    .A3(\adder/adder/_0537_ ),
    .ZN(\adder/adder/_0602_ ));
 NAND2_X1 \adder/adder/_1412_  (.A1(\adder/adder/_0599_ ),
    .A2(\adder/adder/_0602_ ),
    .ZN(\adder/adder/_0603_ ));
 NAND2_X1 \adder/adder/_1413_  (.A1(\adder/adder/_0566_ ),
    .A2(\adder/adder/_0452_ ),
    .ZN(\adder/adder/_0604_ ));
 NAND2_X1 \adder/adder/_1414_  (.A1(\adder/adder/_0577_ ),
    .A2(\adder/adder/_0451_ ),
    .ZN(\adder/adder/_0605_ ));
 NAND2_X1 \adder/adder/_1415_  (.A1(\adder/adder/_0604_ ),
    .A2(\adder/adder/_0605_ ),
    .ZN(\adder/adder/_0606_ ));
 NAND3_X1 \adder/adder/_1416_  (.A1(\adder/adder/_0596_ ),
    .A2(\adder/adder/_0603_ ),
    .A3(\adder/adder/_0606_ ),
    .ZN(\adder/adder/_0607_ ));
 OAI21_X1 \adder/adder/_1417_  (.A(\adder/adder/_0501_ ),
    .B1(\adder/adder/_0593_ ),
    .B2(\adder/adder/_0607_ ),
    .ZN(\adder/adder/_0608_ ));
 NAND2_X1 \adder/adder/_1418_  (.A1(\adder/adder/_0588_ ),
    .A2(\adder/adder/_0452_ ),
    .ZN(\adder/adder/_0609_ ));
 NAND2_X1 \adder/adder/_1419_  (.A1(net245),
    .A2(\operand_fp16_fp32[19] ),
    .ZN(\adder/adder/_0610_ ));
 OAI21_X1 \adder/adder/_1420_  (.A(\adder/adder/_0610_ ),
    .B1(\adder/adder/_0322_ ),
    .B2(net242),
    .ZN(\adder/adder/_0611_ ));
 NAND3_X1 \adder/adder/_1421_  (.A1(net255),
    .A2(\adder/adder/_0611_ ),
    .A3(\adder/adder/_0511_ ),
    .ZN(\adder/adder/_0612_ ));
 NAND2_X1 \adder/adder/_1422_  (.A1(\adder/adder/_0612_ ),
    .A2(\adder/adder/_0451_ ),
    .ZN(\adder/adder/_0613_ ));
 NAND2_X1 \adder/adder/_1423_  (.A1(\adder/adder/_0609_ ),
    .A2(\adder/adder/_0613_ ),
    .ZN(\adder/adder/_0614_ ));
 NAND3_X1 \adder/adder/_1424_  (.A1(\adder/adder/_0614_ ),
    .A2(\adder/adder/_0569_ ),
    .A3(\adder/adder/_0572_ ),
    .ZN(\adder/adder/_0615_ ));
 NAND2_X1 \adder/adder/_1425_  (.A1(\adder/adder/_0615_ ),
    .A2(\adder/adder/_0537_ ),
    .ZN(\adder/adder/_0616_ ));
 NAND2_X1 \adder/adder/_1426_  (.A1(net245),
    .A2(\adder/adder/_0309_ ),
    .ZN(\adder/adder/_0617_ ));
 OAI21_X1 \adder/adder/_1427_  (.A(\adder/adder/_0617_ ),
    .B1(net30),
    .B2(net245),
    .ZN(\adder/adder/_0618_ ));
 INV_X1 \adder/adder/_1428_  (.A(\adder/adder/_0618_ ),
    .ZN(\adder/adder/_0619_ ));
 NAND3_X1 \adder/adder/_1429_  (.A1(net255),
    .A2(\adder/adder/_0619_ ),
    .A3(\adder/adder/_0511_ ),
    .ZN(\adder/adder/_0620_ ));
 NAND2_X1 \adder/adder/_1430_  (.A1(\adder/adder/_0620_ ),
    .A2(\adder/adder/_0452_ ),
    .ZN(\adder/adder/_0621_ ));
 NAND2_X1 \adder/adder/_1431_  (.A1(net242),
    .A2(\operand_fp16_fp32[22] ),
    .ZN(\adder/adder/_0622_ ));
 OAI21_X2 \adder/adder/_1432_  (.A(\adder/adder/_0622_ ),
    .B1(\adder/adder/_0302_ ),
    .B2(net242),
    .ZN(\adder/adder/_0623_ ));
 NAND3_X1 \adder/adder/_1433_  (.A1(net255),
    .A2(\adder/adder/_0623_ ),
    .A3(\adder/adder/_0511_ ),
    .ZN(\adder/adder/_0624_ ));
 NAND2_X1 \adder/adder/_1434_  (.A1(\adder/adder/_0624_ ),
    .A2(\adder/adder/_0451_ ),
    .ZN(\adder/adder/_0625_ ));
 NAND2_X1 \adder/adder/_1435_  (.A1(\adder/adder/_0621_ ),
    .A2(\adder/adder/_0625_ ),
    .ZN(\adder/adder/_0626_ ));
 NAND2_X1 \adder/adder/_1436_  (.A1(\adder/adder/_0624_ ),
    .A2(\adder/adder/_0452_ ),
    .ZN(\adder/adder/_0627_ ));
 NAND2_X1 \adder/adder/_1437_  (.A1(\adder/adder/_0414_ ),
    .A2(\adder/adder/_0338_ ),
    .ZN(\adder/adder/_0628_ ));
 OAI21_X1 \adder/adder/_1438_  (.A(\adder/adder/_0628_ ),
    .B1(\adder/hb_a_d ),
    .B2(\adder/adder/_0414_ ),
    .ZN(\adder/adder/_0629_ ));
 INV_X1 \adder/adder/_1439_  (.A(\adder/adder/_0629_ ),
    .ZN(\adder/adder/_0630_ ));
 NAND3_X1 \adder/adder/_1440_  (.A1(net255),
    .A2(\adder/adder/_0630_ ),
    .A3(\adder/adder/_0511_ ),
    .ZN(\adder/adder/_0631_ ));
 NAND2_X1 \adder/adder/_1441_  (.A1(\adder/adder/_0631_ ),
    .A2(\adder/adder/_0451_ ),
    .ZN(\adder/adder/_0632_ ));
 NAND2_X1 \adder/adder/_1442_  (.A1(\adder/adder/_0627_ ),
    .A2(\adder/adder/_0632_ ),
    .ZN(\adder/adder/_0633_ ));
 NAND3_X1 \adder/adder/_1443_  (.A1(\adder/adder/_0626_ ),
    .A2(\adder/adder/_0633_ ),
    .A3(\adder/adder/_0584_ ),
    .ZN(\adder/adder/_0634_ ));
 NAND2_X1 \adder/adder/_1444_  (.A1(\adder/adder/_0634_ ),
    .A2(\adder/adder/_0538_ ),
    .ZN(\adder/adder/_0635_ ));
 AND2_X4 \adder/adder/_1445_  (.A1(\adder/adder/_0506_ ),
    .A2(\adder/adder/_0511_ ),
    .ZN(\adder/adder/_0636_ ));
 BUF_X1 output57 (.A(net57),
    .Z(result_o[17]));
 NAND2_X1 \adder/adder/_1447_  (.A1(net251),
    .A2(\adder/adder/_0313_ ),
    .ZN(\adder/adder/_0638_ ));
 OAI21_X1 \adder/adder/_1448_  (.A(\adder/adder/_0638_ ),
    .B1(net29),
    .B2(net251),
    .ZN(\adder/adder/_0639_ ));
 INV_X1 \adder/adder/_1449_  (.A(\adder/adder/_0639_ ),
    .ZN(\adder/adder/_0640_ ));
 NAND2_X1 \adder/adder/_1450_  (.A1(\adder/adder/_0636_ ),
    .A2(\adder/adder/_0640_ ),
    .ZN(\adder/adder/_0641_ ));
 NAND2_X1 \adder/adder/_1451_  (.A1(\adder/adder/_0641_ ),
    .A2(\adder/adder/_0452_ ),
    .ZN(\adder/adder/_0642_ ));
 NAND2_X1 \adder/adder/_1452_  (.A1(\adder/adder/_0620_ ),
    .A2(\adder/adder/_0451_ ),
    .ZN(\adder/adder/_0643_ ));
 NAND2_X1 \adder/adder/_1453_  (.A1(\adder/adder/_0642_ ),
    .A2(\adder/adder/_0643_ ),
    .ZN(\adder/adder/_0644_ ));
 NAND2_X1 \adder/adder/_1454_  (.A1(\adder/adder/_0641_ ),
    .A2(\adder/adder/_0451_ ),
    .ZN(\adder/adder/_0645_ ));
 NAND2_X1 \adder/adder/_1455_  (.A1(\adder/adder/_0612_ ),
    .A2(\adder/adder/_0452_ ),
    .ZN(\adder/adder/_0646_ ));
 NAND2_X1 \adder/adder/_1456_  (.A1(\adder/adder/_0645_ ),
    .A2(\adder/adder/_0646_ ),
    .ZN(\adder/adder/_0647_ ));
 NAND2_X1 \adder/adder/_1457_  (.A1(\adder/adder/_0644_ ),
    .A2(\adder/adder/_0647_ ),
    .ZN(\adder/adder/_0648_ ));
 NAND2_X1 \adder/adder/_1458_  (.A1(\adder/adder/_0590_ ),
    .A2(\adder/adder/_0606_ ),
    .ZN(\adder/adder/_0649_ ));
 NOR2_X1 \adder/adder/_1459_  (.A1(\adder/adder/_0648_ ),
    .A2(\adder/adder/_0649_ ),
    .ZN(\adder/adder/_0650_ ));
 NAND3_X1 \adder/adder/_1460_  (.A1(\adder/adder/_0616_ ),
    .A2(\adder/adder/_0635_ ),
    .A3(\adder/adder/_0650_ ),
    .ZN(\adder/adder/_0651_ ));
 INV_X1 \adder/adder/_1461_  (.A(\adder/adder/_0501_ ),
    .ZN(\adder/adder/_0652_ ));
 NAND2_X1 \adder/adder/_1462_  (.A1(\adder/adder/_0651_ ),
    .A2(\adder/adder/_0652_ ),
    .ZN(\adder/adder/_0653_ ));
 MUX2_X1 \adder/adder/_1463_  (.A(\adder/adder/_0584_ ),
    .B(\adder/adder/_0614_ ),
    .S(\adder/adder/_0538_ ),
    .Z(\adder/adder/_0654_ ));
 NAND3_X1 \adder/adder/_1464_  (.A1(\adder/adder/_0608_ ),
    .A2(\adder/adder/_0653_ ),
    .A3(\adder/adder/_0654_ ),
    .ZN(\adder/adder/_0655_ ));
 XNOR2_X1 \adder/adder/_1465_  (.A(\adder/adder/_0500_ ),
    .B(\adder/adder/_0421_ ),
    .ZN(\adder/adder/_0656_ ));
 INV_X1 \adder/adder/_1466_  (.A(\adder/adder/_0656_ ),
    .ZN(\adder/adder/_0657_ ));
 NAND2_X1 \adder/adder/_1467_  (.A1(\adder/adder/_0655_ ),
    .A2(\adder/adder/_0657_ ),
    .ZN(\adder/adder/_0658_ ));
 NAND2_X1 \adder/adder/_1468_  (.A1(net242),
    .A2(\adder/adder/_0244_ ),
    .ZN(\adder/adder/_0659_ ));
 OAI21_X1 \adder/adder/_1469_  (.A(\adder/adder/_0659_ ),
    .B1(net44),
    .B2(net245),
    .ZN(\adder/adder/_0660_ ));
 INV_X1 \adder/adder/_1470_  (.A(\adder/adder/_0660_ ),
    .ZN(\adder/adder/_0661_ ));
 NAND3_X1 \adder/adder/_1471_  (.A1(\adder/adder/_0636_ ),
    .A2(net85),
    .A3(\adder/adder/_0661_ ),
    .ZN(\adder/adder/_0662_ ));
 NAND2_X1 \adder/adder/_1472_  (.A1(net242),
    .A2(\adder/adder/_0218_ ),
    .ZN(\adder/adder/_0663_ ));
 OAI21_X2 \adder/adder/_1473_  (.A(\adder/adder/_0663_ ),
    .B1(net43),
    .B2(net242),
    .ZN(\adder/adder/_0664_ ));
 INV_X1 \adder/adder/_1474_  (.A(\adder/adder/_0664_ ),
    .ZN(\adder/adder/_0665_ ));
 NAND3_X1 \adder/adder/_1475_  (.A1(\adder/adder/_0636_ ),
    .A2(\adder/adder/_0452_ ),
    .A3(\adder/adder/_0665_ ),
    .ZN(\adder/adder/_0666_ ));
 AND2_X1 \adder/adder/_1476_  (.A1(\adder/adder/_0662_ ),
    .A2(\adder/adder/_0666_ ),
    .ZN(\adder/adder/_0667_ ));
 NAND2_X1 \adder/adder/_1477_  (.A1(net239),
    .A2(net204),
    .ZN(\adder/adder/_0668_ ));
 INV_X1 \adder/adder/_1478_  (.A(net42),
    .ZN(\adder/adder/_0669_ ));
 OAI21_X2 \adder/adder/_1479_  (.A(\adder/adder/_0668_ ),
    .B1(\adder/adder/_0669_ ),
    .B2(net242),
    .ZN(\adder/adder/_0670_ ));
 NAND2_X1 \adder/adder/_1480_  (.A1(\adder/adder/_0636_ ),
    .A2(\adder/adder/_0670_ ),
    .ZN(\adder/adder/_0671_ ));
 NAND2_X1 \adder/adder/_1481_  (.A1(\adder/adder/_0671_ ),
    .A2(\adder/adder/_0452_ ),
    .ZN(\adder/adder/_0672_ ));
 NAND2_X1 \adder/adder/_1482_  (.A1(\adder/adder/_0636_ ),
    .A2(\adder/adder/_0665_ ),
    .ZN(\adder/adder/_0673_ ));
 NAND2_X1 \adder/adder/_1483_  (.A1(\adder/adder/_0673_ ),
    .A2(net85),
    .ZN(\adder/adder/_0674_ ));
 NAND2_X1 \adder/adder/_1484_  (.A1(\adder/adder/_0672_ ),
    .A2(\adder/adder/_0674_ ),
    .ZN(\adder/adder/_0675_ ));
 NAND3_X1 \adder/adder/_1485_  (.A1(\adder/adder/_0667_ ),
    .A2(\adder/adder/_0675_ ),
    .A3(\adder/adder/_0538_ ),
    .ZN(\adder/adder/_0676_ ));
 NAND3_X1 \adder/adder/_1486_  (.A1(\adder/adder/_0636_ ),
    .A2(net85),
    .A3(\adder/adder/_0670_ ),
    .ZN(\adder/adder/_0677_ ));
 NAND2_X1 \adder/adder/_1487_  (.A1(net242),
    .A2(\adder/adder/_0138_ ),
    .ZN(\adder/adder/_0678_ ));
 OAI21_X2 \adder/adder/_1488_  (.A(\adder/adder/_0678_ ),
    .B1(net28),
    .B2(net242),
    .ZN(\adder/adder/_0679_ ));
 INV_X1 \adder/adder/_1489_  (.A(\adder/adder/_0679_ ),
    .ZN(\adder/adder/_0680_ ));
 NAND4_X1 \adder/adder/_1490_  (.A1(net255),
    .A2(\adder/adder/_0452_ ),
    .A3(\adder/adder/_0680_ ),
    .A4(\adder/adder/_0511_ ),
    .ZN(\adder/adder/_0681_ ));
 NAND2_X1 \adder/adder/_1491_  (.A1(\adder/adder/_0414_ ),
    .A2(\adder/adder/_0116_ ),
    .ZN(\adder/adder/_0682_ ));
 OAI21_X1 \adder/adder/_1492_  (.A(\adder/adder/_0682_ ),
    .B1(net205),
    .B2(\adder/adder/_0414_ ),
    .ZN(\adder/adder/_0683_ ));
 INV_X1 \adder/adder/_1493_  (.A(\adder/adder/_0683_ ),
    .ZN(\adder/adder/_0684_ ));
 NAND2_X1 \adder/adder/_1494_  (.A1(\adder/adder/_0636_ ),
    .A2(\adder/adder/_0684_ ),
    .ZN(\adder/adder/_0685_ ));
 NAND4_X1 \adder/adder/_1495_  (.A1(\adder/adder/_0677_ ),
    .A2(\adder/adder/_0537_ ),
    .A3(\adder/adder/_0681_ ),
    .A4(\adder/adder/_0685_ ),
    .ZN(\adder/adder/_0686_ ));
 NAND3_X1 \adder/adder/_1496_  (.A1(\adder/adder/_0676_ ),
    .A2(\adder/adder/_0652_ ),
    .A3(\adder/adder/_0686_ ),
    .ZN(\adder/adder/_0687_ ));
 NAND2_X1 \adder/adder/_1497_  (.A1(net242),
    .A2(\adder/adder/_0149_ ),
    .ZN(\adder/adder/_0688_ ));
 OAI21_X1 \adder/adder/_1498_  (.A(\adder/adder/_0688_ ),
    .B1(net17),
    .B2(net242),
    .ZN(\adder/adder/_0689_ ));
 OAI21_X1 \adder/adder/_1499_  (.A(\adder/adder/_0689_ ),
    .B1(\adder/adder/_0679_ ),
    .B2(\adder/adder/_0452_ ),
    .ZN(\adder/adder/_0690_ ));
 NAND2_X1 \adder/adder/_1500_  (.A1(\adder/adder/_0636_ ),
    .A2(\adder/adder/_0690_ ),
    .ZN(\adder/adder/_0691_ ));
 NOR2_X1 \adder/adder/_1501_  (.A1(\adder/adder/_0691_ ),
    .A2(\adder/adder/_0537_ ),
    .ZN(\adder/adder/_0692_ ));
 NAND2_X1 \adder/adder/_1502_  (.A1(\adder/adder/_0692_ ),
    .A2(\adder/adder/_0501_ ),
    .ZN(\adder/adder/_0693_ ));
 NAND2_X1 \adder/adder/_1503_  (.A1(\adder/adder/_0687_ ),
    .A2(\adder/adder/_0693_ ),
    .ZN(\adder/adder/_0694_ ));
 INV_X1 \adder/adder/_1504_  (.A(\adder/adder/_0694_ ),
    .ZN(\adder/adder/_0695_ ));
 NAND2_X1 \adder/adder/_1505_  (.A1(\adder/adder/_0676_ ),
    .A2(\adder/adder/_0686_ ),
    .ZN(\adder/adder/_0696_ ));
 NAND2_X1 \adder/adder/_1506_  (.A1(\adder/adder/_0691_ ),
    .A2(\adder/adder/_0537_ ),
    .ZN(\adder/adder/_0697_ ));
 NAND3_X1 \adder/adder/_1507_  (.A1(\adder/adder/_0677_ ),
    .A2(\adder/adder/_0685_ ),
    .A3(\adder/adder/_0681_ ),
    .ZN(\adder/adder/_0698_ ));
 OAI21_X2 \adder/adder/_1508_  (.A(\adder/adder/_0697_ ),
    .B1(\adder/adder/_0698_ ),
    .B2(\adder/adder/_0537_ ),
    .ZN(\adder/adder/_0699_ ));
 NAND2_X1 \adder/adder/_1509_  (.A1(\adder/adder/_0696_ ),
    .A2(\adder/adder/_0699_ ),
    .ZN(\adder/adder/_0700_ ));
 NAND2_X1 \adder/adder/_1510_  (.A1(\adder/adder/_0700_ ),
    .A2(\adder/adder/_0501_ ),
    .ZN(\adder/adder/_0701_ ));
 NAND3_X1 \adder/adder/_1511_  (.A1(\adder/adder/_0636_ ),
    .A2(\adder/adder/_0452_ ),
    .A3(\adder/adder/_0661_ ),
    .ZN(\adder/adder/_0702_ ));
 NAND2_X1 \adder/adder/_1512_  (.A1(\adder/adder/_0414_ ),
    .A2(\adder/adder/_0072_ ),
    .ZN(\adder/adder/_0703_ ));
 OAI21_X1 \adder/adder/_1513_  (.A(\adder/adder/_0703_ ),
    .B1(net206),
    .B2(\adder/adder/_0414_ ),
    .ZN(\adder/adder/_0704_ ));
 INV_X1 \adder/adder/_1514_  (.A(\adder/adder/_0704_ ),
    .ZN(\adder/adder/_0705_ ));
 NAND2_X1 \adder/adder/_1515_  (.A1(\adder/adder/_0636_ ),
    .A2(\adder/adder/_0705_ ),
    .ZN(\adder/adder/_0706_ ));
 NAND2_X1 \adder/adder/_1516_  (.A1(net251),
    .A2(\adder/adder/_0050_ ),
    .ZN(\adder/adder/_0707_ ));
 OAI21_X1 \adder/adder/_1517_  (.A(\adder/adder/_0707_ ),
    .B1(net46),
    .B2(net245),
    .ZN(\adder/adder/_0708_ ));
 INV_X1 \adder/adder/_1518_  (.A(\adder/adder/_0708_ ),
    .ZN(\adder/adder/_0709_ ));
 NAND2_X1 \adder/adder/_1519_  (.A1(\adder/adder/_0636_ ),
    .A2(\adder/adder/_0709_ ),
    .ZN(\adder/adder/_0710_ ));
 OAI211_X2 \adder/adder/_1520_  (.A(\adder/adder/_0702_ ),
    .B(\adder/adder/_0706_ ),
    .C1(\adder/adder/_0452_ ),
    .C2(\adder/adder/_0710_ ),
    .ZN(\adder/adder/_0711_ ));
 NAND3_X1 \adder/adder/_1521_  (.A1(\adder/adder/_0667_ ),
    .A2(\adder/adder/_0675_ ),
    .A3(\adder/adder/_0537_ ),
    .ZN(\adder/adder/_0712_ ));
 NAND2_X1 \adder/adder/_1522_  (.A1(\adder/adder/_0710_ ),
    .A2(\adder/adder/_0452_ ),
    .ZN(\adder/adder/_0713_ ));
 NAND2_X1 \adder/adder/_1523_  (.A1(net251),
    .A2(\adder/adder/_0276_ ),
    .ZN(\adder/adder/_0714_ ));
 OAI21_X1 \adder/adder/_1524_  (.A(\adder/adder/_0714_ ),
    .B1(net47),
    .B2(net245),
    .ZN(\adder/adder/_0715_ ));
 INV_X1 \adder/adder/_1525_  (.A(\adder/adder/_0715_ ),
    .ZN(\adder/adder/_0716_ ));
 NAND2_X1 \adder/adder/_1526_  (.A1(\adder/adder/_0636_ ),
    .A2(\adder/adder/_0716_ ),
    .ZN(\adder/adder/_0717_ ));
 NAND2_X1 \adder/adder/_1527_  (.A1(\adder/adder/_0717_ ),
    .A2(net85),
    .ZN(\adder/adder/_0718_ ));
 NAND2_X1 \adder/adder/_1528_  (.A1(\adder/adder/_0713_ ),
    .A2(\adder/adder/_0718_ ),
    .ZN(\adder/adder/_0719_ ));
 NAND2_X1 \adder/adder/_1529_  (.A1(\adder/adder/_0717_ ),
    .A2(\adder/adder/_0452_ ),
    .ZN(\adder/adder/_0720_ ));
 NAND2_X1 \adder/adder/_1530_  (.A1(\adder/adder/_0550_ ),
    .A2(net85),
    .ZN(\adder/adder/_0721_ ));
 NAND2_X1 \adder/adder/_1531_  (.A1(\adder/adder/_0720_ ),
    .A2(\adder/adder/_0721_ ),
    .ZN(\adder/adder/_0722_ ));
 NAND3_X1 \adder/adder/_1532_  (.A1(\adder/adder/_0719_ ),
    .A2(\adder/adder/_0722_ ),
    .A3(\adder/adder/_0538_ ),
    .ZN(\adder/adder/_0723_ ));
 AOI21_X1 \adder/adder/_1533_  (.A(\adder/adder/_0711_ ),
    .B1(\adder/adder/_0712_ ),
    .B2(\adder/adder/_0723_ ),
    .ZN(\adder/adder/_0724_ ));
 NAND3_X1 \adder/adder/_1534_  (.A1(\adder/adder/_0695_ ),
    .A2(\adder/adder/_0701_ ),
    .A3(\adder/adder/_0724_ ),
    .ZN(\adder/adder/_0725_ ));
 NAND3_X1 \adder/adder/_1535_  (.A1(\adder/adder/_0719_ ),
    .A2(\adder/adder/_0722_ ),
    .A3(\adder/adder/_0537_ ),
    .ZN(\adder/adder/_0726_ ));
 NAND3_X1 \adder/adder/_1536_  (.A1(\adder/adder/_0546_ ),
    .A2(\adder/adder/_0553_ ),
    .A3(\adder/adder/_0538_ ),
    .ZN(\adder/adder/_0727_ ));
 NAND2_X1 \adder/adder/_1537_  (.A1(\adder/adder/_0726_ ),
    .A2(\adder/adder/_0727_ ),
    .ZN(\adder/adder/_0728_ ));
 INV_X1 \adder/adder/_1538_  (.A(\adder/adder/_0692_ ),
    .ZN(\adder/adder/_0729_ ));
 NAND3_X1 \adder/adder/_1539_  (.A1(\adder/adder/_0728_ ),
    .A2(\adder/adder/_0556_ ),
    .A3(\adder/adder/_0729_ ),
    .ZN(\adder/adder/_0730_ ));
 NAND2_X1 \adder/adder/_1540_  (.A1(\adder/adder/_0730_ ),
    .A2(\adder/adder/_0652_ ),
    .ZN(\adder/adder/_0731_ ));
 AOI21_X1 \adder/adder/_1541_  (.A(\adder/adder/_0501_ ),
    .B1(\adder/adder/_0599_ ),
    .B2(\adder/adder/_0602_ ),
    .ZN(\adder/adder/_0732_ ));
 NAND3_X1 \adder/adder/_1542_  (.A1(\adder/adder/_0699_ ),
    .A2(\adder/adder/_0732_ ),
    .A3(\adder/adder/_0596_ ),
    .ZN(\adder/adder/_0733_ ));
 NAND2_X1 \adder/adder/_1543_  (.A1(\adder/adder/_0728_ ),
    .A2(\adder/adder/_0501_ ),
    .ZN(\adder/adder/_0734_ ));
 NAND2_X1 \adder/adder/_1544_  (.A1(\adder/adder/_0733_ ),
    .A2(\adder/adder/_0734_ ),
    .ZN(\adder/adder/_0735_ ));
 NAND2_X1 \adder/adder/_1545_  (.A1(\adder/adder/_0731_ ),
    .A2(\adder/adder/_0735_ ),
    .ZN(\adder/adder/_0736_ ));
 NOR2_X1 \adder/adder/_1546_  (.A1(\adder/adder/_0725_ ),
    .A2(\adder/adder/_0736_ ),
    .ZN(\adder/adder/_0737_ ));
 NAND2_X1 \adder/adder/_1547_  (.A1(\adder/adder/_0658_ ),
    .A2(\adder/adder/_0737_ ),
    .ZN(\adder/adder/_0738_ ));
 INV_X1 \adder/adder/_1548_  (.A(\adder/adder/_0442_ ),
    .ZN(\adder/adder/_0739_ ));
 INV_X1 \adder/adder/_1549_  (.A(\adder/adder/_0500_ ),
    .ZN(\adder/adder/_0740_ ));
 BUF_X1 output56 (.A(net56),
    .Z(result_o[16]));
 OAI21_X1 \adder/adder/_1551_  (.A(\adder/adder/_0739_ ),
    .B1(\adder/adder/_0740_ ),
    .B2(net265),
    .ZN(\adder/adder/_0742_ ));
 NAND2_X1 \adder/adder/_1552_  (.A1(\adder/adder/_0742_ ),
    .A2(\adder/adder/_0502_ ),
    .ZN(\adder/adder/_0743_ ));
 INV_X1 \adder/adder/_1553_  (.A(\adder/adder/_0743_ ),
    .ZN(\adder/adder/_0744_ ));
 NAND2_X1 \adder/adder/_1554_  (.A1(\adder/adder/_0738_ ),
    .A2(\adder/adder/_0744_ ),
    .ZN(\adder/adder/_0745_ ));
 NAND2_X1 \adder/adder/_1555_  (.A1(\adder/adder/_0743_ ),
    .A2(\adder/adder/_0657_ ),
    .ZN(\adder/adder/_0746_ ));
 NAND2_X1 \adder/adder/_1556_  (.A1(\adder/adder/_0695_ ),
    .A2(\adder/adder/_0699_ ),
    .ZN(\adder/adder/_0747_ ));
 INV_X1 \adder/adder/_1557_  (.A(\adder/adder/_0747_ ),
    .ZN(\adder/adder/_0748_ ));
 OAI21_X1 \adder/adder/_1558_  (.A(\adder/adder/_0712_ ),
    .B1(\adder/adder/_0711_ ),
    .B2(\adder/adder/_0537_ ),
    .ZN(\adder/adder/_0749_ ));
 INV_X1 \adder/adder/_1559_  (.A(\adder/adder/_0749_ ),
    .ZN(\adder/adder/_0750_ ));
 OAI21_X1 \adder/adder/_1560_  (.A(\adder/adder/_0652_ ),
    .B1(\adder/adder/_0750_ ),
    .B2(\adder/adder/_0692_ ),
    .ZN(\adder/adder/_0751_ ));
 AOI21_X1 \adder/adder/_1561_  (.A(\adder/adder/_0746_ ),
    .B1(\adder/adder/_0748_ ),
    .B2(\adder/adder/_0751_ ),
    .ZN(\adder/adder/_0752_ ));
 NOR2_X4 \adder/adder/_1562_  (.A1(\adder/adder/_0437_ ),
    .A2(\adder/adder/_0739_ ),
    .ZN(\adder/adder/_0753_ ));
 BUF_X1 output55 (.A(net55),
    .Z(result_o[15]));
 BUF_X1 output54 (.A(net54),
    .Z(result_o[14]));
 BUF_X1 output53 (.A(net53),
    .Z(result_o[13]));
 BUF_X1 output52 (.A(net52),
    .Z(result_o[12]));
 BUF_X1 output51 (.A(net51),
    .Z(result_o[11]));
 NOR2_X1 \adder/adder/_1568_  (.A1(\adder/adder/_0498_ ),
    .A2(net267),
    .ZN(\adder/adder/_0759_ ));
 NAND4_X1 \adder/adder/_1569_  (.A1(\adder/adder/_0753_ ),
    .A2(\adder/adder/_0421_ ),
    .A3(net85),
    .A4(\adder/adder/_0759_ ),
    .ZN(\adder/adder/_0760_ ));
 INV_X8 \adder/adder/_1570_  (.A(\adder/adder/_0474_ ),
    .ZN(\adder/adder/_0761_ ));
 BUF_X1 output50 (.A(net50),
    .Z(result_o[10]));
 NAND4_X2 \adder/adder/_1572_  (.A1(\adder/adder/_0760_ ),
    .A2(\adder/adder/_0761_ ),
    .A3(\adder/adder/_0436_ ),
    .A4(\adder/adder/_0502_ ),
    .ZN(\adder/adder/_0763_ ));
 NOR2_X1 \adder/adder/_1573_  (.A1(\adder/adder/_0752_ ),
    .A2(\adder/adder/_0763_ ),
    .ZN(\adder/adder/_0764_ ));
 NAND2_X1 \adder/adder/_1574_  (.A1(\adder/adder/_0745_ ),
    .A2(\adder/adder/_0764_ ),
    .ZN(\adder/adder/_0765_ ));
 NAND2_X4 \adder/adder/_1575_  (.A1(\adder/adder/_0477_ ),
    .A2(\adder/adder/_0495_ ),
    .ZN(\adder/adder/_0766_ ));
 INV_X4 \adder/adder/_1576_  (.A(\adder/adder/_0766_ ),
    .ZN(\adder/adder/_0767_ ));
 BUF_X1 output49 (.A(net49),
    .Z(result_o[0]));
 INV_X1 \adder/adder/_1578_  (.A(\adder/adder/_0689_ ),
    .ZN(\adder/adder/_0769_ ));
 NOR4_X1 \adder/adder/_1579_  (.A1(\adder/adder/_0684_ ),
    .A2(\adder/adder/_0680_ ),
    .A3(\adder/adder/_0769_ ),
    .A4(\adder/adder/_0670_ ),
    .ZN(\adder/adder/_0770_ ));
 NOR4_X1 \adder/adder/_1580_  (.A1(\adder/adder/_0665_ ),
    .A2(\adder/adder/_0705_ ),
    .A3(\adder/adder/_0661_ ),
    .A4(\adder/adder/_0709_ ),
    .ZN(\adder/adder/_0771_ ));
 NOR4_X1 \adder/adder/_1581_  (.A1(\adder/adder/_0549_ ),
    .A2(\adder/adder/_0716_ ),
    .A3(\adder/adder/_0542_ ),
    .A4(\adder/adder/_0510_ ),
    .ZN(\adder/adder/_0772_ ));
 NOR4_X1 \adder/adder/_1582_  (.A1(\adder/adder/_0520_ ),
    .A2(\adder/adder/_0531_ ),
    .A3(\adder/adder/_0564_ ),
    .A4(\adder/adder/_0558_ ),
    .ZN(\adder/adder/_0773_ ));
 AND4_X1 \adder/adder/_1583_  (.A1(\adder/adder/_0770_ ),
    .A2(\adder/adder/_0771_ ),
    .A3(\adder/adder/_0772_ ),
    .A4(\adder/adder/_0773_ ),
    .ZN(\adder/adder/_0774_ ));
 NOR4_X1 \adder/adder/_1584_  (.A1(\adder/adder/_0630_ ),
    .A2(\adder/adder/_0640_ ),
    .A3(\adder/adder/_0619_ ),
    .A4(\adder/adder/_0623_ ),
    .ZN(\adder/adder/_0775_ ));
 NOR4_X1 \adder/adder/_1585_  (.A1(\adder/adder/_0581_ ),
    .A2(\adder/adder/_0576_ ),
    .A3(\adder/adder/_0611_ ),
    .A4(\adder/adder/_0587_ ),
    .ZN(\adder/adder/_0776_ ));
 NAND4_X2 \adder/adder/_1586_  (.A1(\adder/adder/_0774_ ),
    .A2(\adder/adder/_0763_ ),
    .A3(\adder/adder/_0775_ ),
    .A4(\adder/adder/_0776_ ),
    .ZN(\adder/adder/_0777_ ));
 NAND3_X1 \adder/adder/_1587_  (.A1(\adder/adder/_0765_ ),
    .A2(\adder/adder/_0767_ ),
    .A3(\adder/adder/_0777_ ),
    .ZN(\adder/adder/_0778_ ));
 OAI21_X1 \adder/adder/_1588_  (.A(net85),
    .B1(\adder/adder/_0474_ ),
    .B2(\adder/adder/_0664_ ),
    .ZN(\adder/adder/_0779_ ));
 NOR2_X1 \adder/adder/_1589_  (.A1(\adder/adder/_0474_ ),
    .A2(\adder/adder/_0660_ ),
    .ZN(\adder/adder/_0780_ ));
 OAI21_X1 \adder/adder/_1590_  (.A(\adder/adder/_0779_ ),
    .B1(net85),
    .B2(\adder/adder/_0780_ ),
    .ZN(\adder/adder/_0781_ ));
 INV_X1 \adder/adder/_1591_  (.A(\adder/adder/_0781_ ),
    .ZN(\adder/adder/_0782_ ));
 BUF_X1 input48 (.A(operand_fp32_i[9]),
    .Z(net48));
 NAND2_X1 \adder/adder/_1593_  (.A1(\adder/adder/_0782_ ),
    .A2(\adder/adder/_0450_ ),
    .ZN(\adder/adder/_0784_ ));
 NAND2_X1 \adder/adder/_1594_  (.A1(\adder/adder/_0761_ ),
    .A2(\adder/adder/_0670_ ),
    .ZN(\adder/adder/_0785_ ));
 NAND2_X1 \adder/adder/_1595_  (.A1(\adder/adder/_0785_ ),
    .A2(\adder/adder/_0452_ ),
    .ZN(\adder/adder/_0786_ ));
 NAND2_X1 \adder/adder/_1596_  (.A1(\adder/adder/_0761_ ),
    .A2(\adder/adder/_0684_ ),
    .ZN(\adder/adder/_0787_ ));
 NAND2_X1 \adder/adder/_1597_  (.A1(\adder/adder/_0787_ ),
    .A2(net85),
    .ZN(\adder/adder/_0788_ ));
 NAND2_X1 \adder/adder/_1598_  (.A1(\adder/adder/_0786_ ),
    .A2(\adder/adder/_0788_ ),
    .ZN(\adder/adder/_0789_ ));
 OAI21_X1 \adder/adder/_1599_  (.A(\adder/adder/_0784_ ),
    .B1(\adder/adder/_0450_ ),
    .B2(\adder/adder/_0789_ ),
    .ZN(\adder/adder/_0790_ ));
 NAND2_X1 \adder/adder/_1600_  (.A1(\adder/adder/_0761_ ),
    .A2(\adder/adder/_0769_ ),
    .ZN(\adder/adder/_0791_ ));
 NAND2_X1 \adder/adder/_1601_  (.A1(\adder/adder/_0791_ ),
    .A2(net85),
    .ZN(\adder/adder/_0792_ ));
 NOR2_X1 \adder/adder/_1602_  (.A1(\adder/adder/_0474_ ),
    .A2(\adder/adder/_0679_ ),
    .ZN(\adder/adder/_0793_ ));
 OAI21_X1 \adder/adder/_1603_  (.A(\adder/adder/_0792_ ),
    .B1(net85),
    .B2(\adder/adder/_0793_ ),
    .ZN(\adder/adder/_0794_ ));
 INV_X1 \adder/adder/_1604_  (.A(\adder/adder/_0794_ ),
    .ZN(\adder/adder/_0795_ ));
 AOI22_X1 \adder/adder/_1605_  (.A1(\adder/adder/_0790_ ),
    .A2(\adder/adder/_0498_ ),
    .B1(\adder/adder/_0795_ ),
    .B2(\adder/adder/_0759_ ),
    .ZN(\adder/adder/_0796_ ));
 NAND2_X1 \adder/adder/_1606_  (.A1(\adder/adder/_0796_ ),
    .A2(net252),
    .ZN(\adder/adder/_0797_ ));
 BUF_X1 input47 (.A(operand_fp32_i[8]),
    .Z(net47));
 NAND2_X1 \adder/adder/_1608_  (.A1(\adder/adder/_0761_ ),
    .A2(\adder/adder/_0709_ ),
    .ZN(\adder/adder/_0799_ ));
 BUF_X1 input46 (.A(operand_fp32_i[7]),
    .Z(net46));
 NAND2_X1 \adder/adder/_1610_  (.A1(\adder/adder/_0799_ ),
    .A2(\adder/adder/_0452_ ),
    .ZN(\adder/adder/_0801_ ));
 NAND2_X1 \adder/adder/_1611_  (.A1(\adder/adder/_0761_ ),
    .A2(\adder/adder/_0705_ ),
    .ZN(\adder/adder/_0802_ ));
 NAND2_X1 \adder/adder/_1612_  (.A1(\adder/adder/_0802_ ),
    .A2(net85),
    .ZN(\adder/adder/_0803_ ));
 BUF_X1 input45 (.A(operand_fp32_i[6]),
    .Z(net45));
 NAND3_X1 \adder/adder/_1614_  (.A1(\adder/adder/_0801_ ),
    .A2(\adder/adder/_0803_ ),
    .A3(\adder/adder/_0449_ ),
    .ZN(\adder/adder/_0805_ ));
 NAND2_X1 \adder/adder/_1615_  (.A1(\adder/adder/_0761_ ),
    .A2(\adder/adder/_0716_ ),
    .ZN(\adder/adder/_0806_ ));
 NAND2_X1 \adder/adder/_1616_  (.A1(\adder/adder/_0806_ ),
    .A2(net85),
    .ZN(\adder/adder/_0807_ ));
 NOR2_X1 \adder/adder/_1617_  (.A1(\adder/adder/_0474_ ),
    .A2(\adder/adder/_0548_ ),
    .ZN(\adder/adder/_0808_ ));
 OAI21_X1 \adder/adder/_1618_  (.A(\adder/adder/_0807_ ),
    .B1(net85),
    .B2(\adder/adder/_0808_ ),
    .ZN(\adder/adder/_0809_ ));
 OAI21_X1 \adder/adder/_1619_  (.A(\adder/adder/_0805_ ),
    .B1(\adder/adder/_0809_ ),
    .B2(\adder/adder/_0449_ ),
    .ZN(\adder/adder/_0810_ ));
 OR2_X1 \adder/adder/_1620_  (.A1(\adder/adder/_0810_ ),
    .A2(\adder/adder/_0498_ ),
    .ZN(\adder/adder/_0811_ ));
 BUF_X1 input44 (.A(operand_fp32_i[5]),
    .Z(net44));
 NAND2_X1 \adder/adder/_1622_  (.A1(\adder/adder/_0761_ ),
    .A2(\adder/adder/_0510_ ),
    .ZN(\adder/adder/_0813_ ));
 NAND2_X1 \adder/adder/_1623_  (.A1(\adder/adder/_0813_ ),
    .A2(\adder/adder/_0452_ ),
    .ZN(\adder/adder/_0814_ ));
 NAND2_X1 \adder/adder/_1624_  (.A1(\adder/adder/_0761_ ),
    .A2(\adder/adder/_0542_ ),
    .ZN(\adder/adder/_0815_ ));
 NAND2_X1 \adder/adder/_1625_  (.A1(\adder/adder/_0815_ ),
    .A2(net85),
    .ZN(\adder/adder/_0816_ ));
 NAND2_X1 \adder/adder/_1626_  (.A1(\adder/adder/_0814_ ),
    .A2(\adder/adder/_0816_ ),
    .ZN(\adder/adder/_0817_ ));
 INV_X1 \adder/adder/_1627_  (.A(\adder/adder/_0817_ ),
    .ZN(\adder/adder/_0818_ ));
 NAND2_X1 \adder/adder/_1628_  (.A1(\adder/adder/_0818_ ),
    .A2(net267),
    .ZN(\adder/adder/_0819_ ));
 NAND2_X1 \adder/adder/_1629_  (.A1(\adder/adder/_0761_ ),
    .A2(\adder/adder/_0531_ ),
    .ZN(\adder/adder/_0820_ ));
 NAND2_X1 \adder/adder/_1630_  (.A1(\adder/adder/_0820_ ),
    .A2(\adder/adder/_0452_ ),
    .ZN(\adder/adder/_0821_ ));
 NOR2_X1 \adder/adder/_1631_  (.A1(\adder/adder/_0474_ ),
    .A2(\adder/adder/_0519_ ),
    .ZN(\adder/adder/_0822_ ));
 OAI21_X1 \adder/adder/_1632_  (.A(\adder/adder/_0821_ ),
    .B1(\adder/adder/_0452_ ),
    .B2(\adder/adder/_0822_ ),
    .ZN(\adder/adder/_0823_ ));
 OAI21_X1 \adder/adder/_1633_  (.A(\adder/adder/_0819_ ),
    .B1(net267),
    .B2(\adder/adder/_0823_ ),
    .ZN(\adder/adder/_0824_ ));
 OAI21_X1 \adder/adder/_1634_  (.A(\adder/adder/_0811_ ),
    .B1(net272),
    .B2(\adder/adder/_0824_ ),
    .ZN(\adder/adder/_0825_ ));
 NAND2_X1 \adder/adder/_1635_  (.A1(\adder/adder/_0825_ ),
    .A2(\adder/adder/_0421_ ),
    .ZN(\adder/adder/_0826_ ));
 BUF_X1 input43 (.A(operand_fp32_i[4]),
    .Z(net43));
 NAND3_X1 \adder/adder/_1637_  (.A1(\adder/adder/_0797_ ),
    .A2(\adder/adder/_0826_ ),
    .A3(net266),
    .ZN(\adder/adder/_0828_ ));
 NAND3_X1 \adder/adder/_1638_  (.A1(\adder/adder/_0761_ ),
    .A2(net85),
    .A3(\adder/adder/_0623_ ),
    .ZN(\adder/adder/_0829_ ));
 NAND2_X1 \adder/adder/_1639_  (.A1(\adder/adder/_0761_ ),
    .A2(\adder/adder/_0630_ ),
    .ZN(\adder/adder/_0830_ ));
 OAI21_X1 \adder/adder/_1640_  (.A(\adder/adder/_0829_ ),
    .B1(net85),
    .B2(\adder/adder/_0830_ ),
    .ZN(\adder/adder/_0831_ ));
 NAND2_X1 \adder/adder/_1641_  (.A1(\adder/adder/_0831_ ),
    .A2(\adder/adder/_0449_ ),
    .ZN(\adder/adder/_0832_ ));
 NOR2_X1 \adder/adder/_1642_  (.A1(\adder/adder/_0832_ ),
    .A2(\adder/adder/_0498_ ),
    .ZN(\adder/adder/_0833_ ));
 NAND2_X1 \adder/adder/_1643_  (.A1(\adder/adder/_0833_ ),
    .A2(\adder/adder/_0421_ ),
    .ZN(\adder/adder/_0834_ ));
 NAND2_X1 \adder/adder/_1644_  (.A1(\adder/adder/_0761_ ),
    .A2(\adder/adder/_0558_ ),
    .ZN(\adder/adder/_0835_ ));
 NAND2_X1 \adder/adder/_1645_  (.A1(\adder/adder/_0835_ ),
    .A2(net85),
    .ZN(\adder/adder/_0836_ ));
 NOR2_X1 \adder/adder/_1646_  (.A1(\adder/adder/_0474_ ),
    .A2(\adder/adder/_0563_ ),
    .ZN(\adder/adder/_0837_ ));
 OAI21_X1 \adder/adder/_1647_  (.A(\adder/adder/_0836_ ),
    .B1(net85),
    .B2(\adder/adder/_0837_ ),
    .ZN(\adder/adder/_0838_ ));
 INV_X2 \adder/adder/_1648_  (.A(\adder/adder/_0838_ ),
    .ZN(\adder/adder/_0839_ ));
 NAND2_X1 \adder/adder/_1649_  (.A1(\adder/adder/_0839_ ),
    .A2(net267),
    .ZN(\adder/adder/_0840_ ));
 NAND3_X1 \adder/adder/_1650_  (.A1(\adder/adder/_0761_ ),
    .A2(net85),
    .A3(\adder/adder/_0576_ ),
    .ZN(\adder/adder/_0841_ ));
 NAND2_X1 \adder/adder/_1651_  (.A1(\adder/adder/_0761_ ),
    .A2(\adder/adder/_0581_ ),
    .ZN(\adder/adder/_0842_ ));
 OAI21_X1 \adder/adder/_1652_  (.A(\adder/adder/_0841_ ),
    .B1(net85),
    .B2(\adder/adder/_0842_ ),
    .ZN(\adder/adder/_0843_ ));
 BUF_X1 input42 (.A(operand_fp32_i[3]),
    .Z(net42));
 NAND2_X1 \adder/adder/_1654_  (.A1(\adder/adder/_0843_ ),
    .A2(\adder/adder/_0450_ ),
    .ZN(\adder/adder/_0845_ ));
 NAND3_X1 \adder/adder/_1655_  (.A1(\adder/adder/_0840_ ),
    .A2(\adder/adder/_0458_ ),
    .A3(\adder/adder/_0845_ ),
    .ZN(\adder/adder/_0846_ ));
 NAND2_X1 \adder/adder/_1656_  (.A1(\adder/adder/_0761_ ),
    .A2(\adder/adder/_0640_ ),
    .ZN(\adder/adder/_0847_ ));
 INV_X1 \adder/adder/_1657_  (.A(\adder/adder/_0847_ ),
    .ZN(\adder/adder/_0848_ ));
 NAND2_X1 \adder/adder/_1658_  (.A1(\adder/adder/_0848_ ),
    .A2(\adder/adder/_0451_ ),
    .ZN(\adder/adder/_0849_ ));
 NAND2_X1 \adder/adder/_1659_  (.A1(\adder/adder/_0761_ ),
    .A2(\adder/adder/_0619_ ),
    .ZN(\adder/adder/_0850_ ));
 OAI21_X1 \adder/adder/_1660_  (.A(\adder/adder/_0849_ ),
    .B1(\adder/adder/_0451_ ),
    .B2(\adder/adder/_0850_ ),
    .ZN(\adder/adder/_0851_ ));
 NAND2_X1 \adder/adder/_1661_  (.A1(\adder/adder/_0851_ ),
    .A2(\adder/adder/_0450_ ),
    .ZN(\adder/adder/_0852_ ));
 NAND3_X1 \adder/adder/_1662_  (.A1(\adder/adder/_0761_ ),
    .A2(net85),
    .A3(\adder/adder/_0587_ ),
    .ZN(\adder/adder/_0853_ ));
 NAND2_X1 \adder/adder/_1663_  (.A1(\adder/adder/_0761_ ),
    .A2(\adder/adder/_0611_ ),
    .ZN(\adder/adder/_0854_ ));
 OAI21_X1 \adder/adder/_1664_  (.A(\adder/adder/_0853_ ),
    .B1(net85),
    .B2(\adder/adder/_0854_ ),
    .ZN(\adder/adder/_0855_ ));
 NAND2_X1 \adder/adder/_1665_  (.A1(\adder/adder/_0855_ ),
    .A2(\adder/adder/_0449_ ),
    .ZN(\adder/adder/_0856_ ));
 NAND2_X1 \adder/adder/_1666_  (.A1(\adder/adder/_0852_ ),
    .A2(\adder/adder/_0856_ ),
    .ZN(\adder/adder/_0857_ ));
 OAI21_X1 \adder/adder/_1667_  (.A(\adder/adder/_0846_ ),
    .B1(net272),
    .B2(\adder/adder/_0857_ ),
    .ZN(\adder/adder/_0858_ ));
 OAI21_X1 \adder/adder/_1668_  (.A(\adder/adder/_0834_ ),
    .B1(\adder/adder/_0858_ ),
    .B2(\adder/adder/_0421_ ),
    .ZN(\adder/adder/_0859_ ));
 NAND2_X1 \adder/adder/_1669_  (.A1(\adder/adder/_0859_ ),
    .A2(\adder/adder/_0753_ ),
    .ZN(\adder/adder/_0860_ ));
 NAND2_X1 \adder/adder/_1670_  (.A1(\adder/adder/_0828_ ),
    .A2(\adder/adder/_0860_ ),
    .ZN(\adder/adder/_0861_ ));
 XNOR2_X1 \adder/adder/_1671_  (.A(\adder/adder/_0861_ ),
    .B(\adder/adder/_0767_ ),
    .ZN(\adder/adder/_0862_ ));
 NOR2_X4 \adder/adder/_1672_  (.A1(\adder/adder/_0494_ ),
    .A2(\adder/adder/_0477_ ),
    .ZN(\adder/adder/_0863_ ));
 INV_X8 \adder/adder/_1673_  (.A(\adder/adder/_0863_ ),
    .ZN(\adder/adder/_0864_ ));
 BUF_X1 input41 (.A(operand_fp32_i[31]),
    .Z(net41));
 BUF_X1 input40 (.A(operand_fp32_i[30]),
    .Z(net40));
 NAND2_X1 \adder/adder/_1676_  (.A1(\adder/adder/_0862_ ),
    .A2(\adder/adder/_0864_ ),
    .ZN(\adder/adder/_0867_ ));
 NAND3_X1 \adder/adder/_1677_  (.A1(\adder/adder/_0761_ ),
    .A2(net85),
    .A3(\adder/adder/_0531_ ),
    .ZN(\adder/adder/_0868_ ));
 OAI21_X1 \adder/adder/_1678_  (.A(\adder/adder/_0868_ ),
    .B1(net85),
    .B2(\adder/adder/_0835_ ),
    .ZN(\adder/adder/_0869_ ));
 NAND2_X1 \adder/adder/_1679_  (.A1(\adder/adder/_0869_ ),
    .A2(\adder/adder/_0450_ ),
    .ZN(\adder/adder/_0870_ ));
 NAND2_X1 \adder/adder/_1680_  (.A1(\adder/adder/_0813_ ),
    .A2(net85),
    .ZN(\adder/adder/_0871_ ));
 OAI21_X1 \adder/adder/_1681_  (.A(\adder/adder/_0871_ ),
    .B1(net85),
    .B2(\adder/adder/_0822_ ),
    .ZN(\adder/adder/_0872_ ));
 OAI21_X1 \adder/adder/_1682_  (.A(\adder/adder/_0870_ ),
    .B1(\adder/adder/_0450_ ),
    .B2(\adder/adder/_0872_ ),
    .ZN(\adder/adder/_0873_ ));
 BUF_X1 input39 (.A(operand_fp32_i[2]),
    .Z(net39));
 OR2_X1 \adder/adder/_1684_  (.A1(\adder/adder/_0873_ ),
    .A2(net272),
    .ZN(\adder/adder/_0875_ ));
 NAND2_X1 \adder/adder/_1685_  (.A1(\adder/adder/_0806_ ),
    .A2(\adder/adder/_0452_ ),
    .ZN(\adder/adder/_0876_ ));
 INV_X1 \adder/adder/_1686_  (.A(\adder/adder/_0799_ ),
    .ZN(\adder/adder/_0877_ ));
 OAI21_X1 \adder/adder/_1687_  (.A(\adder/adder/_0876_ ),
    .B1(\adder/adder/_0452_ ),
    .B2(\adder/adder/_0877_ ),
    .ZN(\adder/adder/_0878_ ));
 OR2_X1 \adder/adder/_1688_  (.A1(\adder/adder/_0878_ ),
    .A2(\adder/adder/_0450_ ),
    .ZN(\adder/adder/_0879_ ));
 NAND2_X1 \adder/adder/_1689_  (.A1(\adder/adder/_0815_ ),
    .A2(\adder/adder/_0452_ ),
    .ZN(\adder/adder/_0880_ ));
 OAI21_X1 \adder/adder/_1690_  (.A(\adder/adder/_0880_ ),
    .B1(\adder/adder/_0452_ ),
    .B2(\adder/adder/_0808_ ),
    .ZN(\adder/adder/_0881_ ));
 OAI21_X1 \adder/adder/_1691_  (.A(\adder/adder/_0879_ ),
    .B1(net267),
    .B2(\adder/adder/_0881_ ),
    .ZN(\adder/adder/_0882_ ));
 OAI21_X1 \adder/adder/_1692_  (.A(\adder/adder/_0875_ ),
    .B1(\adder/adder/_0498_ ),
    .B2(\adder/adder/_0882_ ),
    .ZN(\adder/adder/_0883_ ));
 NAND2_X1 \adder/adder/_1693_  (.A1(\adder/adder/_0883_ ),
    .A2(\adder/adder/_0421_ ),
    .ZN(\adder/adder/_0884_ ));
 OAI21_X1 \adder/adder/_1694_  (.A(net267),
    .B1(\adder/adder/_0791_ ),
    .B2(net85),
    .ZN(\adder/adder/_0885_ ));
 NAND3_X1 \adder/adder/_1695_  (.A1(\adder/adder/_0761_ ),
    .A2(net85),
    .A3(\adder/adder/_0680_ ),
    .ZN(\adder/adder/_0886_ ));
 OAI21_X1 \adder/adder/_1696_  (.A(\adder/adder/_0886_ ),
    .B1(net85),
    .B2(\adder/adder/_0787_ ),
    .ZN(\adder/adder/_0887_ ));
 OAI21_X1 \adder/adder/_1697_  (.A(\adder/adder/_0885_ ),
    .B1(\adder/adder/_0887_ ),
    .B2(net267),
    .ZN(\adder/adder/_0888_ ));
 NAND2_X1 \adder/adder/_1698_  (.A1(\adder/adder/_0888_ ),
    .A2(net254),
    .ZN(\adder/adder/_0889_ ));
 NAND2_X1 \adder/adder/_1699_  (.A1(\adder/adder/_0780_ ),
    .A2(net85),
    .ZN(\adder/adder/_0890_ ));
 OAI21_X1 \adder/adder/_1700_  (.A(\adder/adder/_0890_ ),
    .B1(net85),
    .B2(\adder/adder/_0802_ ),
    .ZN(\adder/adder/_0891_ ));
 NAND2_X1 \adder/adder/_1701_  (.A1(\adder/adder/_0891_ ),
    .A2(\adder/adder/_0450_ ),
    .ZN(\adder/adder/_0892_ ));
 NAND2_X1 \adder/adder/_1702_  (.A1(\adder/adder/_0785_ ),
    .A2(net85),
    .ZN(\adder/adder/_0893_ ));
 OAI21_X1 \adder/adder/_1703_  (.A(\adder/adder/_0452_ ),
    .B1(\adder/adder/_0474_ ),
    .B2(\adder/adder/_0664_ ),
    .ZN(\adder/adder/_0894_ ));
 NAND2_X1 \adder/adder/_1704_  (.A1(\adder/adder/_0893_ ),
    .A2(\adder/adder/_0894_ ),
    .ZN(\adder/adder/_0895_ ));
 OAI21_X1 \adder/adder/_1705_  (.A(\adder/adder/_0892_ ),
    .B1(\adder/adder/_0450_ ),
    .B2(\adder/adder/_0895_ ),
    .ZN(\adder/adder/_0896_ ));
 OAI21_X1 \adder/adder/_1706_  (.A(\adder/adder/_0889_ ),
    .B1(\adder/adder/_0896_ ),
    .B2(net254),
    .ZN(\adder/adder/_0897_ ));
 NAND2_X1 \adder/adder/_1707_  (.A1(\adder/adder/_0897_ ),
    .A2(net265),
    .ZN(\adder/adder/_0898_ ));
 NAND3_X1 \adder/adder/_1708_  (.A1(\adder/adder/_0884_ ),
    .A2(net266),
    .A3(\adder/adder/_0898_ ),
    .ZN(\adder/adder/_0899_ ));
 NOR3_X1 \adder/adder/_1709_  (.A1(\adder/adder/_0830_ ),
    .A2(\adder/adder/_0452_ ),
    .A3(\adder/adder/_0450_ ),
    .ZN(\adder/adder/_0900_ ));
 INV_X1 \adder/adder/_1710_  (.A(\adder/adder/_0900_ ),
    .ZN(\adder/adder/_0901_ ));
 NOR2_X1 \adder/adder/_1711_  (.A1(\adder/adder/_0901_ ),
    .A2(\adder/adder/_0498_ ),
    .ZN(\adder/adder/_0902_ ));
 NAND2_X1 \adder/adder/_1712_  (.A1(\adder/adder/_0902_ ),
    .A2(\adder/adder/_0421_ ),
    .ZN(\adder/adder/_0903_ ));
 NAND2_X1 \adder/adder/_1713_  (.A1(\adder/adder/_0761_ ),
    .A2(\adder/adder/_0623_ ),
    .ZN(\adder/adder/_0904_ ));
 NAND2_X1 \adder/adder/_1714_  (.A1(\adder/adder/_0904_ ),
    .A2(\adder/adder/_0452_ ),
    .ZN(\adder/adder/_0905_ ));
 INV_X1 \adder/adder/_1715_  (.A(\adder/adder/_0850_ ),
    .ZN(\adder/adder/_0906_ ));
 OAI21_X1 \adder/adder/_1716_  (.A(\adder/adder/_0905_ ),
    .B1(\adder/adder/_0452_ ),
    .B2(\adder/adder/_0906_ ),
    .ZN(\adder/adder/_0907_ ));
 INV_X1 \adder/adder/_1717_  (.A(\adder/adder/_0907_ ),
    .ZN(\adder/adder/_0908_ ));
 NAND2_X1 \adder/adder/_1718_  (.A1(\adder/adder/_0908_ ),
    .A2(\adder/adder/_0450_ ),
    .ZN(\adder/adder/_0909_ ));
 NAND2_X1 \adder/adder/_1719_  (.A1(\adder/adder/_0854_ ),
    .A2(net85),
    .ZN(\adder/adder/_0910_ ));
 OAI21_X1 \adder/adder/_1720_  (.A(\adder/adder/_0910_ ),
    .B1(net85),
    .B2(\adder/adder/_0848_ ),
    .ZN(\adder/adder/_0911_ ));
 OAI21_X1 \adder/adder/_1721_  (.A(\adder/adder/_0909_ ),
    .B1(\adder/adder/_0450_ ),
    .B2(\adder/adder/_0911_ ),
    .ZN(\adder/adder/_0912_ ));
 NAND2_X1 \adder/adder/_1722_  (.A1(\adder/adder/_0912_ ),
    .A2(\adder/adder/_0498_ ),
    .ZN(\adder/adder/_0913_ ));
 NAND3_X1 \adder/adder/_1723_  (.A1(\adder/adder/_0761_ ),
    .A2(\adder/adder/_0452_ ),
    .A3(\adder/adder/_0587_ ),
    .ZN(\adder/adder/_0914_ ));
 OAI21_X1 \adder/adder/_1724_  (.A(\adder/adder/_0914_ ),
    .B1(\adder/adder/_0452_ ),
    .B2(\adder/adder/_0842_ ),
    .ZN(\adder/adder/_0915_ ));
 NAND2_X1 \adder/adder/_1725_  (.A1(\adder/adder/_0915_ ),
    .A2(\adder/adder/_0450_ ),
    .ZN(\adder/adder/_0916_ ));
 OAI21_X1 \adder/adder/_1726_  (.A(\adder/adder/_0452_ ),
    .B1(\adder/adder/_0474_ ),
    .B2(\adder/adder/_0575_ ),
    .ZN(\adder/adder/_0917_ ));
 OAI21_X1 \adder/adder/_1727_  (.A(\adder/adder/_0917_ ),
    .B1(\adder/adder/_0452_ ),
    .B2(\adder/adder/_0837_ ),
    .ZN(\adder/adder/_0918_ ));
 OAI21_X1 \adder/adder/_1728_  (.A(\adder/adder/_0916_ ),
    .B1(\adder/adder/_0450_ ),
    .B2(\adder/adder/_0918_ ),
    .ZN(\adder/adder/_0919_ ));
 NAND2_X1 \adder/adder/_1729_  (.A1(\adder/adder/_0919_ ),
    .A2(net254),
    .ZN(\adder/adder/_0920_ ));
 AND2_X1 \adder/adder/_1730_  (.A1(\adder/adder/_0913_ ),
    .A2(\adder/adder/_0920_ ),
    .ZN(\adder/adder/_0921_ ));
 OAI21_X1 \adder/adder/_1731_  (.A(\adder/adder/_0903_ ),
    .B1(\adder/adder/_0921_ ),
    .B2(\adder/adder/_0421_ ),
    .ZN(\adder/adder/_0922_ ));
 NAND2_X1 \adder/adder/_1732_  (.A1(\adder/adder/_0922_ ),
    .A2(\adder/adder/_0753_ ),
    .ZN(\adder/adder/_0923_ ));
 NAND2_X1 \adder/adder/_1733_  (.A1(\adder/adder/_0899_ ),
    .A2(\adder/adder/_0923_ ),
    .ZN(\adder/adder/_0924_ ));
 NAND2_X1 \adder/adder/_1734_  (.A1(\adder/adder/_0924_ ),
    .A2(\adder/adder/_0767_ ),
    .ZN(\adder/adder/_0925_ ));
 NAND3_X1 \adder/adder/_1735_  (.A1(\adder/adder/_0899_ ),
    .A2(\adder/adder/_0923_ ),
    .A3(\adder/adder/_0766_ ),
    .ZN(\adder/adder/_0926_ ));
 AOI21_X2 \adder/adder/_1736_  (.A(\adder/adder/_0863_ ),
    .B1(\adder/adder/_0925_ ),
    .B2(\adder/adder/_0926_ ),
    .ZN(\adder/adder/_0927_ ));
 NAND2_X1 \adder/adder/_1737_  (.A1(\adder/adder/_0801_ ),
    .A2(\adder/adder/_0803_ ),
    .ZN(\adder/adder/_0928_ ));
 NAND2_X1 \adder/adder/_1738_  (.A1(\adder/adder/_0928_ ),
    .A2(\adder/adder/_0450_ ),
    .ZN(\adder/adder/_0929_ ));
 OAI21_X1 \adder/adder/_1739_  (.A(\adder/adder/_0929_ ),
    .B1(\adder/adder/_0782_ ),
    .B2(\adder/adder/_0450_ ),
    .ZN(\adder/adder/_0930_ ));
 AND2_X1 \adder/adder/_1740_  (.A1(\adder/adder/_0930_ ),
    .A2(\adder/adder/_0498_ ),
    .ZN(\adder/adder/_0931_ ));
 NAND2_X1 \adder/adder/_1741_  (.A1(\adder/adder/_0794_ ),
    .A2(net267),
    .ZN(\adder/adder/_0932_ ));
 NAND2_X1 \adder/adder/_1742_  (.A1(\adder/adder/_0789_ ),
    .A2(\adder/adder/_0450_ ),
    .ZN(\adder/adder/_0933_ ));
 AOI21_X1 \adder/adder/_1743_  (.A(\adder/adder/_0498_ ),
    .B1(\adder/adder/_0932_ ),
    .B2(\adder/adder/_0933_ ),
    .ZN(\adder/adder/_0934_ ));
 OAI21_X1 \adder/adder/_1744_  (.A(net265),
    .B1(\adder/adder/_0931_ ),
    .B2(\adder/adder/_0934_ ),
    .ZN(\adder/adder/_0935_ ));
 NAND2_X1 \adder/adder/_1745_  (.A1(\adder/adder/_0823_ ),
    .A2(\adder/adder/_0449_ ),
    .ZN(\adder/adder/_0936_ ));
 OAI21_X1 \adder/adder/_1746_  (.A(\adder/adder/_0936_ ),
    .B1(net267),
    .B2(\adder/adder/_0839_ ),
    .ZN(\adder/adder/_0937_ ));
 NAND2_X1 \adder/adder/_1747_  (.A1(\adder/adder/_0937_ ),
    .A2(\adder/adder/_0498_ ),
    .ZN(\adder/adder/_0938_ ));
 NAND2_X1 \adder/adder/_1748_  (.A1(\adder/adder/_0809_ ),
    .A2(\adder/adder/_0449_ ),
    .ZN(\adder/adder/_0939_ ));
 OAI21_X1 \adder/adder/_1749_  (.A(\adder/adder/_0939_ ),
    .B1(\adder/adder/_0449_ ),
    .B2(\adder/adder/_0818_ ),
    .ZN(\adder/adder/_0940_ ));
 NAND2_X1 \adder/adder/_1750_  (.A1(\adder/adder/_0940_ ),
    .A2(net272),
    .ZN(\adder/adder/_0941_ ));
 NAND2_X1 \adder/adder/_1751_  (.A1(\adder/adder/_0938_ ),
    .A2(\adder/adder/_0941_ ),
    .ZN(\adder/adder/_0942_ ));
 NAND2_X1 \adder/adder/_1752_  (.A1(\adder/adder/_0942_ ),
    .A2(\adder/adder/_0421_ ),
    .ZN(\adder/adder/_0943_ ));
 NAND3_X1 \adder/adder/_1753_  (.A1(\adder/adder/_0935_ ),
    .A2(\adder/adder/_0943_ ),
    .A3(net266),
    .ZN(\adder/adder/_0944_ ));
 MUX2_X1 \adder/adder/_1754_  (.A(\adder/adder/_0831_ ),
    .B(\adder/adder/_0851_ ),
    .S(\adder/adder/_0449_ ),
    .Z(\adder/adder/_0945_ ));
 NAND2_X1 \adder/adder/_1755_  (.A1(\adder/adder/_0945_ ),
    .A2(\adder/adder/_0498_ ),
    .ZN(\adder/adder/_0946_ ));
 MUX2_X1 \adder/adder/_1756_  (.A(\adder/adder/_0843_ ),
    .B(\adder/adder/_0855_ ),
    .S(\adder/adder/_0450_ ),
    .Z(\adder/adder/_0947_ ));
 NAND2_X1 \adder/adder/_1757_  (.A1(\adder/adder/_0947_ ),
    .A2(net254),
    .ZN(\adder/adder/_0948_ ));
 AOI21_X2 \adder/adder/_1758_  (.A(\adder/adder/_0421_ ),
    .B1(\adder/adder/_0946_ ),
    .B2(\adder/adder/_0948_ ),
    .ZN(\adder/adder/_0949_ ));
 NAND2_X1 \adder/adder/_1759_  (.A1(\adder/adder/_0949_ ),
    .A2(\adder/adder/_0753_ ),
    .ZN(\adder/adder/_0950_ ));
 NAND2_X1 \adder/adder/_1760_  (.A1(\adder/adder/_0944_ ),
    .A2(\adder/adder/_0950_ ),
    .ZN(\adder/adder/_0951_ ));
 NAND2_X1 \adder/adder/_1761_  (.A1(\adder/adder/_0951_ ),
    .A2(\adder/adder/_0767_ ),
    .ZN(\adder/adder/_0952_ ));
 NAND3_X1 \adder/adder/_1762_  (.A1(\adder/adder/_0944_ ),
    .A2(\adder/adder/_0950_ ),
    .A3(\adder/adder/_0766_ ),
    .ZN(\adder/adder/_0953_ ));
 NAND2_X1 \adder/adder/_1763_  (.A1(\adder/adder/_0952_ ),
    .A2(\adder/adder/_0953_ ),
    .ZN(\adder/adder/_0954_ ));
 BUF_X1 input38 (.A(operand_fp32_i[29]),
    .Z(net38));
 NAND2_X1 \adder/adder/_1765_  (.A1(\adder/adder/_0414_ ),
    .A2(\adder/adder/_0149_ ),
    .ZN(\adder/adder/_0956_ ));
 OAI21_X1 \adder/adder/_1766_  (.A(\adder/adder/_0956_ ),
    .B1(net17),
    .B2(\adder/adder/_0414_ ),
    .ZN(\adder/adder/_0957_ ));
 XNOR2_X1 \adder/adder/_1767_  (.A(\adder/adder/_0863_ ),
    .B(\adder/adder/_0957_ ),
    .ZN(\adder/adder/_0958_ ));
 INV_X1 \adder/adder/_1768_  (.A(\adder/adder/_0958_ ),
    .ZN(\adder/adder/_0959_ ));
 NAND2_X1 \adder/adder/_1769_  (.A1(\adder/adder/_0954_ ),
    .A2(\adder/adder/_0959_ ),
    .ZN(\adder/adder/_0960_ ));
 NAND3_X1 \adder/adder/_1770_  (.A1(\adder/adder/_0952_ ),
    .A2(\adder/adder/_0953_ ),
    .A3(\adder/adder/_0958_ ),
    .ZN(\adder/adder/_0961_ ));
 NAND2_X1 \adder/adder/_1771_  (.A1(\adder/adder/_0960_ ),
    .A2(\adder/adder/_0961_ ),
    .ZN(\adder/adder/_0962_ ));
 NOR2_X1 \adder/adder/_1772_  (.A1(\adder/adder/_0927_ ),
    .A2(\adder/adder/_0962_ ),
    .ZN(\adder/adder/_0963_ ));
 NAND4_X1 \adder/adder/_1773_  (.A1(\adder/adder/_0778_ ),
    .A2(\adder/adder/_0495_ ),
    .A3(\adder/adder/_0867_ ),
    .A4(\adder/adder/_0963_ ),
    .ZN(\adder/adder/_0964_ ));
 NAND2_X2 \adder/adder/_1774_  (.A1(\adder/adder/_0964_ ),
    .A2(\adder/adder/_0961_ ),
    .ZN(\adder/adder/_0965_ ));
 OR2_X1 \adder/adder/_1775_  (.A1(\adder/adder/_0919_ ),
    .A2(net272),
    .ZN(\adder/adder/_0966_ ));
 OAI21_X1 \adder/adder/_1776_  (.A(\adder/adder/_0966_ ),
    .B1(\adder/adder/_0873_ ),
    .B2(\adder/adder/_0498_ ),
    .ZN(\adder/adder/_0967_ ));
 NAND2_X1 \adder/adder/_1777_  (.A1(\adder/adder/_0967_ ),
    .A2(\adder/adder/_0421_ ),
    .ZN(\adder/adder/_0968_ ));
 NOR2_X1 \adder/adder/_1778_  (.A1(\adder/adder/_0882_ ),
    .A2(net254),
    .ZN(\adder/adder/_0969_ ));
 NOR2_X1 \adder/adder/_1779_  (.A1(\adder/adder/_0896_ ),
    .A2(\adder/adder/_0498_ ),
    .ZN(\adder/adder/_0970_ ));
 OAI21_X1 \adder/adder/_1780_  (.A(net265),
    .B1(\adder/adder/_0969_ ),
    .B2(\adder/adder/_0970_ ),
    .ZN(\adder/adder/_0971_ ));
 NAND3_X1 \adder/adder/_1781_  (.A1(\adder/adder/_0968_ ),
    .A2(\adder/adder/_0971_ ),
    .A3(\adder/adder/_0443_ ),
    .ZN(\adder/adder/_0972_ ));
 NOR2_X1 \adder/adder/_1782_  (.A1(\adder/adder/_0901_ ),
    .A2(net254),
    .ZN(\adder/adder/_0973_ ));
 AOI21_X1 \adder/adder/_1783_  (.A(\adder/adder/_0973_ ),
    .B1(\adder/adder/_0912_ ),
    .B2(net254),
    .ZN(\adder/adder/_0974_ ));
 INV_X1 \adder/adder/_1784_  (.A(\adder/adder/_0974_ ),
    .ZN(\adder/adder/_0975_ ));
 NAND3_X1 \adder/adder/_1785_  (.A1(\adder/adder/_0975_ ),
    .A2(net252),
    .A3(\adder/adder/_0753_ ),
    .ZN(\adder/adder/_0976_ ));
 NAND2_X1 \adder/adder/_1786_  (.A1(\adder/adder/_0972_ ),
    .A2(\adder/adder/_0976_ ),
    .ZN(\adder/adder/_0977_ ));
 XNOR2_X2 \adder/adder/_1787_  (.A(\adder/adder/_0977_ ),
    .B(\adder/adder/_0767_ ),
    .ZN(\adder/adder/_0978_ ));
 NAND2_X1 \adder/adder/_1788_  (.A1(net239),
    .A2(\adder/adder/_0669_ ),
    .ZN(\adder/adder/_0979_ ));
 OAI21_X1 \adder/adder/_1789_  (.A(\adder/adder/_0979_ ),
    .B1(net207),
    .B2(net239),
    .ZN(\adder/adder/_0980_ ));
 XNOR2_X2 \adder/adder/_1790_  (.A(\adder/adder/_0864_ ),
    .B(\adder/adder/_0980_ ),
    .ZN(\adder/adder/_0981_ ));
 XNOR2_X2 \adder/adder/_1791_  (.A(\adder/adder/_0978_ ),
    .B(\adder/adder/_0981_ ),
    .ZN(\adder/adder/_0982_ ));
 MUX2_X1 \adder/adder/_1792_  (.A(\adder/adder/_0930_ ),
    .B(\adder/adder/_0940_ ),
    .S(\adder/adder/_0498_ ),
    .Z(\adder/adder/_0983_ ));
 NAND2_X1 \adder/adder/_1793_  (.A1(\adder/adder/_0983_ ),
    .A2(net265),
    .ZN(\adder/adder/_0984_ ));
 NAND2_X1 \adder/adder/_1794_  (.A1(\adder/adder/_0937_ ),
    .A2(\adder/adder/_0458_ ),
    .ZN(\adder/adder/_0985_ ));
 OAI21_X1 \adder/adder/_1795_  (.A(\adder/adder/_0985_ ),
    .B1(net254),
    .B2(\adder/adder/_0947_ ),
    .ZN(\adder/adder/_0986_ ));
 NAND2_X1 \adder/adder/_1796_  (.A1(\adder/adder/_0986_ ),
    .A2(\adder/adder/_0421_ ),
    .ZN(\adder/adder/_0987_ ));
 NAND3_X1 \adder/adder/_1797_  (.A1(\adder/adder/_0984_ ),
    .A2(net266),
    .A3(\adder/adder/_0987_ ),
    .ZN(\adder/adder/_0988_ ));
 NAND2_X1 \adder/adder/_1798_  (.A1(\adder/adder/_0945_ ),
    .A2(net254),
    .ZN(\adder/adder/_0989_ ));
 INV_X1 \adder/adder/_1799_  (.A(\adder/adder/_0989_ ),
    .ZN(\adder/adder/_0990_ ));
 NAND3_X1 \adder/adder/_1800_  (.A1(\adder/adder/_0990_ ),
    .A2(net265),
    .A3(\adder/adder/_0753_ ),
    .ZN(\adder/adder/_0991_ ));
 NAND2_X1 \adder/adder/_1801_  (.A1(\adder/adder/_0988_ ),
    .A2(\adder/adder/_0991_ ),
    .ZN(\adder/adder/_0992_ ));
 XNOR2_X1 \adder/adder/_1802_  (.A(\adder/adder/_0992_ ),
    .B(\adder/adder/_0767_ ),
    .ZN(\adder/adder/_0993_ ));
 NAND2_X1 \adder/adder/_1803_  (.A1(net242),
    .A2(\adder/adder/_0235_ ),
    .ZN(\adder/adder/_0994_ ));
 OAI21_X1 \adder/adder/_1804_  (.A(\adder/adder/_0994_ ),
    .B1(net208),
    .B2(net239),
    .ZN(\adder/adder/_0995_ ));
 XNOR2_X1 \adder/adder/_1805_  (.A(\adder/adder/_0864_ ),
    .B(\adder/adder/_0995_ ),
    .ZN(\adder/adder/_0996_ ));
 NOR2_X1 \adder/adder/_1806_  (.A1(\adder/adder/_0993_ ),
    .A2(\adder/adder/_0996_ ),
    .ZN(\adder/adder/_0997_ ));
 INV_X1 \adder/adder/_1807_  (.A(\adder/adder/_0997_ ),
    .ZN(\adder/adder/_0998_ ));
 NAND2_X1 \adder/adder/_1808_  (.A1(\adder/adder/_0993_ ),
    .A2(\adder/adder/_0996_ ),
    .ZN(\adder/adder/_0999_ ));
 NAND2_X1 \adder/adder/_1809_  (.A1(\adder/adder/_0998_ ),
    .A2(\adder/adder/_0999_ ),
    .ZN(\adder/adder/_1000_ ));
 NOR2_X1 \adder/adder/_1810_  (.A1(\adder/adder/_0982_ ),
    .A2(\adder/adder/_1000_ ),
    .ZN(\adder/adder/_1001_ ));
 MUX2_X1 \adder/adder/_1811_  (.A(\adder/adder/_0872_ ),
    .B(\adder/adder/_0881_ ),
    .S(\adder/adder/_0449_ ),
    .Z(\adder/adder/_1002_ ));
 NAND2_X1 \adder/adder/_1812_  (.A1(\adder/adder/_1002_ ),
    .A2(\adder/adder/_0458_ ),
    .ZN(\adder/adder/_1003_ ));
 NAND2_X1 \adder/adder/_1813_  (.A1(\adder/adder/_0869_ ),
    .A2(net267),
    .ZN(\adder/adder/_1004_ ));
 OAI21_X1 \adder/adder/_1814_  (.A(\adder/adder/_1004_ ),
    .B1(net267),
    .B2(\adder/adder/_0918_ ),
    .ZN(\adder/adder/_1005_ ));
 OAI21_X1 \adder/adder/_1815_  (.A(\adder/adder/_1003_ ),
    .B1(\adder/adder/_1005_ ),
    .B2(net272),
    .ZN(\adder/adder/_1006_ ));
 NAND2_X1 \adder/adder/_1816_  (.A1(\adder/adder/_1006_ ),
    .A2(\adder/adder/_0421_ ),
    .ZN(\adder/adder/_1007_ ));
 NAND2_X1 \adder/adder/_1817_  (.A1(\adder/adder/_0895_ ),
    .A2(\adder/adder/_0450_ ),
    .ZN(\adder/adder/_1008_ ));
 OAI21_X1 \adder/adder/_1818_  (.A(\adder/adder/_1008_ ),
    .B1(\adder/adder/_0887_ ),
    .B2(\adder/adder/_0450_ ),
    .ZN(\adder/adder/_1009_ ));
 NAND2_X1 \adder/adder/_1819_  (.A1(\adder/adder/_1009_ ),
    .A2(net254),
    .ZN(\adder/adder/_1010_ ));
 NAND2_X1 \adder/adder/_1820_  (.A1(\adder/adder/_0891_ ),
    .A2(net267),
    .ZN(\adder/adder/_1011_ ));
 OAI21_X1 \adder/adder/_1821_  (.A(\adder/adder/_1011_ ),
    .B1(net267),
    .B2(\adder/adder/_0878_ ),
    .ZN(\adder/adder/_1012_ ));
 OAI21_X1 \adder/adder/_1822_  (.A(\adder/adder/_1010_ ),
    .B1(\adder/adder/_1012_ ),
    .B2(net254),
    .ZN(\adder/adder/_1013_ ));
 NAND2_X1 \adder/adder/_1823_  (.A1(\adder/adder/_1013_ ),
    .A2(net265),
    .ZN(\adder/adder/_1014_ ));
 NAND3_X1 \adder/adder/_1824_  (.A1(\adder/adder/_1007_ ),
    .A2(net266),
    .A3(\adder/adder/_1014_ ),
    .ZN(\adder/adder/_1015_ ));
 INV_X1 \adder/adder/_1825_  (.A(\adder/adder/_0830_ ),
    .ZN(\adder/adder/_1016_ ));
 AOI21_X1 \adder/adder/_1826_  (.A(\adder/adder/_0449_ ),
    .B1(\adder/adder/_1016_ ),
    .B2(net85),
    .ZN(\adder/adder/_1017_ ));
 AOI21_X1 \adder/adder/_1827_  (.A(\adder/adder/_1017_ ),
    .B1(\adder/adder/_0907_ ),
    .B2(\adder/adder/_0449_ ),
    .ZN(\adder/adder/_1018_ ));
 NAND2_X1 \adder/adder/_1828_  (.A1(\adder/adder/_0915_ ),
    .A2(\adder/adder/_0449_ ),
    .ZN(\adder/adder/_1019_ ));
 OAI21_X1 \adder/adder/_1829_  (.A(\adder/adder/_1019_ ),
    .B1(\adder/adder/_0449_ ),
    .B2(\adder/adder/_0911_ ),
    .ZN(\adder/adder/_1020_ ));
 MUX2_X1 \adder/adder/_1830_  (.A(\adder/adder/_1018_ ),
    .B(\adder/adder/_1020_ ),
    .S(\adder/adder/_0458_ ),
    .Z(\adder/adder/_1021_ ));
 NAND3_X1 \adder/adder/_1831_  (.A1(\adder/adder/_1021_ ),
    .A2(net265),
    .A3(\adder/adder/_0753_ ),
    .ZN(\adder/adder/_1022_ ));
 NAND2_X1 \adder/adder/_1832_  (.A1(\adder/adder/_1015_ ),
    .A2(\adder/adder/_1022_ ),
    .ZN(\adder/adder/_1023_ ));
 NAND2_X1 \adder/adder/_1833_  (.A1(\adder/adder/_1023_ ),
    .A2(\adder/adder/_0767_ ),
    .ZN(\adder/adder/_1024_ ));
 NAND3_X1 \adder/adder/_1834_  (.A1(\adder/adder/_1015_ ),
    .A2(\adder/adder/_0766_ ),
    .A3(\adder/adder/_1022_ ),
    .ZN(\adder/adder/_1025_ ));
 NAND2_X1 \adder/adder/_1835_  (.A1(\adder/adder/_1024_ ),
    .A2(\adder/adder/_1025_ ),
    .ZN(\adder/adder/_1026_ ));
 NAND2_X1 \adder/adder/_1836_  (.A1(net242),
    .A2(\adder/adder/_0171_ ),
    .ZN(\adder/adder/_1027_ ));
 OAI21_X1 \adder/adder/_1837_  (.A(\adder/adder/_1027_ ),
    .B1(net209),
    .B2(net242),
    .ZN(\adder/adder/_1028_ ));
 XNOR2_X1 \adder/adder/_1838_  (.A(\adder/adder/_0864_ ),
    .B(\adder/adder/_1028_ ),
    .ZN(\adder/adder/_1029_ ));
 OR2_X1 \adder/adder/_1839_  (.A1(\adder/adder/_1026_ ),
    .A2(\adder/adder/_1029_ ),
    .ZN(\adder/adder/_1030_ ));
 NAND2_X1 \adder/adder/_1840_  (.A1(\adder/adder/_1026_ ),
    .A2(\adder/adder/_1029_ ),
    .ZN(\adder/adder/_1031_ ));
 NAND2_X1 \adder/adder/_1841_  (.A1(\adder/adder/_1030_ ),
    .A2(\adder/adder/_1031_ ),
    .ZN(\adder/adder/_1032_ ));
 NOR2_X1 \adder/adder/_1842_  (.A1(\adder/adder/_0790_ ),
    .A2(\adder/adder/_0498_ ),
    .ZN(\adder/adder/_1033_ ));
 NOR2_X1 \adder/adder/_1843_  (.A1(\adder/adder/_0810_ ),
    .A2(net254),
    .ZN(\adder/adder/_1034_ ));
 OAI21_X1 \adder/adder/_1844_  (.A(net265),
    .B1(\adder/adder/_1033_ ),
    .B2(\adder/adder/_1034_ ),
    .ZN(\adder/adder/_1035_ ));
 NAND3_X1 \adder/adder/_1845_  (.A1(\adder/adder/_0840_ ),
    .A2(\adder/adder/_0498_ ),
    .A3(\adder/adder/_0845_ ),
    .ZN(\adder/adder/_1036_ ));
 OAI21_X1 \adder/adder/_1846_  (.A(\adder/adder/_1036_ ),
    .B1(\adder/adder/_0498_ ),
    .B2(\adder/adder/_0824_ ),
    .ZN(\adder/adder/_1037_ ));
 NAND2_X1 \adder/adder/_1847_  (.A1(\adder/adder/_1037_ ),
    .A2(\adder/adder/_0421_ ),
    .ZN(\adder/adder/_1038_ ));
 NAND3_X1 \adder/adder/_1848_  (.A1(\adder/adder/_1035_ ),
    .A2(net266),
    .A3(\adder/adder/_1038_ ),
    .ZN(\adder/adder/_1039_ ));
 NAND2_X1 \adder/adder/_1849_  (.A1(\adder/adder/_0832_ ),
    .A2(\adder/adder/_0498_ ),
    .ZN(\adder/adder/_1040_ ));
 OAI21_X1 \adder/adder/_1850_  (.A(\adder/adder/_1040_ ),
    .B1(\adder/adder/_0857_ ),
    .B2(\adder/adder/_0498_ ),
    .ZN(\adder/adder/_1041_ ));
 OR2_X1 \adder/adder/_1851_  (.A1(\adder/adder/_1041_ ),
    .A2(\adder/adder/_0421_ ),
    .ZN(\adder/adder/_1042_ ));
 INV_X1 \adder/adder/_1852_  (.A(\adder/adder/_1042_ ),
    .ZN(\adder/adder/_1043_ ));
 NAND2_X1 \adder/adder/_1853_  (.A1(\adder/adder/_1043_ ),
    .A2(\adder/adder/_0753_ ),
    .ZN(\adder/adder/_1044_ ));
 NAND2_X1 \adder/adder/_1854_  (.A1(\adder/adder/_1039_ ),
    .A2(\adder/adder/_1044_ ),
    .ZN(\adder/adder/_1045_ ));
 XNOR2_X2 \adder/adder/_1855_  (.A(\adder/adder/_1045_ ),
    .B(\adder/adder/_0767_ ),
    .ZN(\adder/adder/_1046_ ));
 NAND2_X1 \adder/adder/_1856_  (.A1(net239),
    .A2(\adder/adder/_0116_ ),
    .ZN(\adder/adder/_1047_ ));
 OAI21_X1 \adder/adder/_1857_  (.A(\adder/adder/_1047_ ),
    .B1(net210),
    .B2(net242),
    .ZN(\adder/adder/_1048_ ));
 XNOR2_X2 \adder/adder/_1858_  (.A(\adder/adder/_0864_ ),
    .B(\adder/adder/_1048_ ),
    .ZN(\adder/adder/_1049_ ));
 XNOR2_X2 \adder/adder/_1859_  (.A(\adder/adder/_1046_ ),
    .B(\adder/adder/_1049_ ),
    .ZN(\adder/adder/_1050_ ));
 NOR2_X1 \adder/adder/_1860_  (.A1(\adder/adder/_1032_ ),
    .A2(\adder/adder/_1050_ ),
    .ZN(\adder/adder/_1051_ ));
 AND2_X1 \adder/adder/_1861_  (.A1(\adder/adder/_1001_ ),
    .A2(\adder/adder/_1051_ ),
    .ZN(\adder/adder/_1052_ ));
 NAND2_X1 \adder/adder/_1862_  (.A1(\adder/adder/_0965_ ),
    .A2(\adder/adder/_1052_ ),
    .ZN(\adder/adder/_1053_ ));
 NOR2_X1 \adder/adder/_1863_  (.A1(\adder/adder/_0978_ ),
    .A2(\adder/adder/_0981_ ),
    .ZN(\adder/adder/_1054_ ));
 AOI21_X1 \adder/adder/_1864_  (.A(\adder/adder/_0997_ ),
    .B1(\adder/adder/_1054_ ),
    .B2(\adder/adder/_0999_ ),
    .ZN(\adder/adder/_1055_ ));
 INV_X1 \adder/adder/_1865_  (.A(\adder/adder/_1001_ ),
    .ZN(\adder/adder/_1056_ ));
 NOR2_X1 \adder/adder/_1866_  (.A1(\adder/adder/_1046_ ),
    .A2(\adder/adder/_1049_ ),
    .ZN(\adder/adder/_1057_ ));
 INV_X1 \adder/adder/_1867_  (.A(\adder/adder/_1057_ ),
    .ZN(\adder/adder/_1058_ ));
 OAI21_X1 \adder/adder/_1868_  (.A(\adder/adder/_1058_ ),
    .B1(\adder/adder/_1050_ ),
    .B2(\adder/adder/_1030_ ),
    .ZN(\adder/adder/_1059_ ));
 INV_X2 \adder/adder/_1869_  (.A(\adder/adder/_1059_ ),
    .ZN(\adder/adder/_1060_ ));
 OAI21_X1 \adder/adder/_1870_  (.A(\adder/adder/_1055_ ),
    .B1(\adder/adder/_1056_ ),
    .B2(\adder/adder/_1060_ ),
    .ZN(\adder/adder/_1061_ ));
 INV_X2 \adder/adder/_1871_  (.A(\adder/adder/_1061_ ),
    .ZN(\adder/adder/_1062_ ));
 NAND2_X2 \adder/adder/_1872_  (.A1(\adder/adder/_1053_ ),
    .A2(\adder/adder/_1062_ ),
    .ZN(\adder/adder/_1063_ ));
 NAND2_X1 \adder/adder/_1873_  (.A1(\adder/adder/_1002_ ),
    .A2(\adder/adder/_0498_ ),
    .ZN(\adder/adder/_1064_ ));
 OAI21_X1 \adder/adder/_1874_  (.A(\adder/adder/_1064_ ),
    .B1(\adder/adder/_1012_ ),
    .B2(\adder/adder/_0498_ ),
    .ZN(\adder/adder/_1065_ ));
 BUF_X1 input37 (.A(operand_fp32_i[28]),
    .Z(net37));
 NAND2_X1 \adder/adder/_1876_  (.A1(\adder/adder/_1065_ ),
    .A2(net252),
    .ZN(\adder/adder/_1067_ ));
 OR2_X1 \adder/adder/_1877_  (.A1(\adder/adder/_1020_ ),
    .A2(net272),
    .ZN(\adder/adder/_1068_ ));
 OAI21_X1 \adder/adder/_1878_  (.A(\adder/adder/_1068_ ),
    .B1(\adder/adder/_1005_ ),
    .B2(\adder/adder/_0498_ ),
    .ZN(\adder/adder/_1069_ ));
 NAND2_X1 \adder/adder/_1879_  (.A1(\adder/adder/_1069_ ),
    .A2(\adder/adder/_0421_ ),
    .ZN(\adder/adder/_1070_ ));
 NAND3_X1 \adder/adder/_1880_  (.A1(\adder/adder/_1067_ ),
    .A2(\adder/adder/_1070_ ),
    .A3(net253),
    .ZN(\adder/adder/_1071_ ));
 INV_X1 \adder/adder/_1881_  (.A(\adder/adder/_0753_ ),
    .ZN(\adder/adder/_1072_ ));
 NAND2_X1 \adder/adder/_1882_  (.A1(\adder/adder/_1018_ ),
    .A2(net254),
    .ZN(\adder/adder/_1073_ ));
 NOR2_X1 \adder/adder/_1883_  (.A1(\adder/adder/_1073_ ),
    .A2(\adder/adder/_0421_ ),
    .ZN(\adder/adder/_1074_ ));
 INV_X1 \adder/adder/_1884_  (.A(\adder/adder/_1074_ ),
    .ZN(\adder/adder/_1075_ ));
 OAI21_X1 \adder/adder/_1885_  (.A(\adder/adder/_1071_ ),
    .B1(\adder/adder/_1072_ ),
    .B2(\adder/adder/_1075_ ),
    .ZN(\adder/adder/_1076_ ));
 XNOR2_X2 \adder/adder/_1886_  (.A(\adder/adder/_1076_ ),
    .B(\adder/adder/_0767_ ),
    .ZN(\adder/adder/_1077_ ));
 NAND2_X1 \adder/adder/_1887_  (.A1(net239),
    .A2(\adder/adder/_0241_ ),
    .ZN(\adder/adder/_1078_ ));
 OAI21_X1 \adder/adder/_1888_  (.A(\adder/adder/_1078_ ),
    .B1(net211),
    .B2(net239),
    .ZN(\adder/adder/_1079_ ));
 XNOR2_X2 \adder/adder/_1889_  (.A(\adder/adder/_0864_ ),
    .B(\adder/adder/_1079_ ),
    .ZN(\adder/adder/_1080_ ));
 XNOR2_X2 \adder/adder/_1890_  (.A(\adder/adder/_1077_ ),
    .B(\adder/adder/_1080_ ),
    .ZN(\adder/adder/_1081_ ));
 NAND2_X1 \adder/adder/_1891_  (.A1(\adder/adder/_0825_ ),
    .A2(net265),
    .ZN(\adder/adder/_1082_ ));
 NAND2_X1 \adder/adder/_1892_  (.A1(\adder/adder/_0858_ ),
    .A2(\adder/adder/_0421_ ),
    .ZN(\adder/adder/_1083_ ));
 NAND3_X1 \adder/adder/_1893_  (.A1(\adder/adder/_1082_ ),
    .A2(\adder/adder/_1083_ ),
    .A3(net266),
    .ZN(\adder/adder/_1084_ ));
 NAND3_X1 \adder/adder/_1894_  (.A1(\adder/adder/_0833_ ),
    .A2(net265),
    .A3(\adder/adder/_0753_ ),
    .ZN(\adder/adder/_1085_ ));
 NAND2_X1 \adder/adder/_1895_  (.A1(\adder/adder/_1084_ ),
    .A2(\adder/adder/_1085_ ),
    .ZN(\adder/adder/_1086_ ));
 XNOR2_X1 \adder/adder/_1896_  (.A(\adder/adder/_1086_ ),
    .B(\adder/adder/_0767_ ),
    .ZN(\adder/adder/_1087_ ));
 NAND2_X1 \adder/adder/_1897_  (.A1(net239),
    .A2(\adder/adder/_0072_ ),
    .ZN(\adder/adder/_1088_ ));
 OAI21_X1 \adder/adder/_1898_  (.A(\adder/adder/_1088_ ),
    .B1(net212),
    .B2(net242),
    .ZN(\adder/adder/_1089_ ));
 XNOR2_X1 \adder/adder/_1899_  (.A(\adder/adder/_0864_ ),
    .B(\adder/adder/_1089_ ),
    .ZN(\adder/adder/_1090_ ));
 AND2_X1 \adder/adder/_1900_  (.A1(\adder/adder/_1087_ ),
    .A2(\adder/adder/_1090_ ),
    .ZN(\adder/adder/_1091_ ));
 NOR2_X1 \adder/adder/_1901_  (.A1(\adder/adder/_1087_ ),
    .A2(\adder/adder/_1090_ ),
    .ZN(\adder/adder/_1092_ ));
 OR2_X1 \adder/adder/_1902_  (.A1(\adder/adder/_1091_ ),
    .A2(\adder/adder/_1092_ ),
    .ZN(\adder/adder/_1093_ ));
 NOR2_X1 \adder/adder/_1903_  (.A1(\adder/adder/_1081_ ),
    .A2(\adder/adder/_1093_ ),
    .ZN(\adder/adder/_1094_ ));
 NAND2_X1 \adder/adder/_1904_  (.A1(\adder/adder/_0883_ ),
    .A2(net265),
    .ZN(\adder/adder/_1095_ ));
 NAND2_X1 \adder/adder/_1905_  (.A1(\adder/adder/_0921_ ),
    .A2(\adder/adder/_0421_ ),
    .ZN(\adder/adder/_1096_ ));
 NAND3_X1 \adder/adder/_1906_  (.A1(\adder/adder/_1095_ ),
    .A2(\adder/adder/_1096_ ),
    .A3(\adder/adder/_0443_ ),
    .ZN(\adder/adder/_1097_ ));
 INV_X1 \adder/adder/_1907_  (.A(\adder/adder/_0902_ ),
    .ZN(\adder/adder/_1098_ ));
 NOR2_X1 \adder/adder/_1908_  (.A1(\adder/adder/_1098_ ),
    .A2(\adder/adder/_0421_ ),
    .ZN(\adder/adder/_1099_ ));
 INV_X1 \adder/adder/_1909_  (.A(\adder/adder/_1099_ ),
    .ZN(\adder/adder/_1100_ ));
 OAI21_X1 \adder/adder/_1910_  (.A(\adder/adder/_1097_ ),
    .B1(\adder/adder/_1100_ ),
    .B2(\adder/adder/_1072_ ),
    .ZN(\adder/adder/_1101_ ));
 XNOR2_X1 \adder/adder/_1911_  (.A(\adder/adder/_1101_ ),
    .B(\adder/adder/_0767_ ),
    .ZN(\adder/adder/_1102_ ));
 NAND2_X1 \adder/adder/_1912_  (.A1(\adder/adder/_0414_ ),
    .A2(\adder/adder/_0050_ ),
    .ZN(\adder/adder/_1103_ ));
 OAI21_X1 \adder/adder/_1913_  (.A(\adder/adder/_1103_ ),
    .B1(net46),
    .B2(\adder/adder/_0414_ ),
    .ZN(\adder/adder/_1104_ ));
 XNOR2_X2 \adder/adder/_1914_  (.A(\adder/adder/_0864_ ),
    .B(\adder/adder/_1104_ ),
    .ZN(\adder/adder/_1105_ ));
 XNOR2_X2 \adder/adder/_1915_  (.A(\adder/adder/_1102_ ),
    .B(\adder/adder/_1105_ ),
    .ZN(\adder/adder/_1106_ ));
 NAND3_X1 \adder/adder/_1916_  (.A1(\adder/adder/_0946_ ),
    .A2(\adder/adder/_0421_ ),
    .A3(\adder/adder/_0948_ ),
    .ZN(\adder/adder/_0000_ ));
 NAND2_X1 \adder/adder/_1917_  (.A1(\adder/adder/_0942_ ),
    .A2(net252),
    .ZN(\adder/adder/_0001_ ));
 NAND3_X1 \adder/adder/_1918_  (.A1(\adder/adder/_0000_ ),
    .A2(net266),
    .A3(\adder/adder/_0001_ ),
    .ZN(\adder/adder/_0002_ ));
 XNOR2_X2 \adder/adder/_1919_  (.A(\adder/adder/_0002_ ),
    .B(\adder/adder/_0766_ ),
    .ZN(\adder/adder/_0003_ ));
 NAND2_X1 \adder/adder/_1920_  (.A1(net239),
    .A2(\adder/adder/_0278_ ),
    .ZN(\adder/adder/_0004_ ));
 OAI21_X1 \adder/adder/_1921_  (.A(\adder/adder/_0004_ ),
    .B1(net213),
    .B2(net239),
    .ZN(\adder/adder/_0005_ ));
 XNOR2_X2 \adder/adder/_1922_  (.A(\adder/adder/_0864_ ),
    .B(\adder/adder/_0005_ ),
    .ZN(\adder/adder/_0006_ ));
 XNOR2_X2 \adder/adder/_1923_  (.A(\adder/adder/_0003_ ),
    .B(\adder/adder/_0006_ ),
    .ZN(\adder/adder/_0007_ ));
 NOR2_X1 \adder/adder/_1924_  (.A1(\adder/adder/_1106_ ),
    .A2(\adder/adder/_0007_ ),
    .ZN(\adder/adder/_0008_ ));
 NAND2_X1 \adder/adder/_1925_  (.A1(\adder/adder/_1094_ ),
    .A2(\adder/adder/_0008_ ),
    .ZN(\adder/adder/_0009_ ));
 NAND2_X1 \adder/adder/_1926_  (.A1(\adder/adder/_1021_ ),
    .A2(\adder/adder/_0421_ ),
    .ZN(\adder/adder/_0010_ ));
 OAI21_X1 \adder/adder/_1927_  (.A(\adder/adder/_0010_ ),
    .B1(\adder/adder/_0421_ ),
    .B2(\adder/adder/_1006_ ),
    .ZN(\adder/adder/_0011_ ));
 NAND2_X1 \adder/adder/_1928_  (.A1(\adder/adder/_0011_ ),
    .A2(net253),
    .ZN(\adder/adder/_0012_ ));
 XNOR2_X1 \adder/adder/_1929_  (.A(\adder/adder/_0012_ ),
    .B(\adder/adder/_0766_ ),
    .ZN(\adder/adder/_0013_ ));
 NAND2_X1 \adder/adder/_1930_  (.A1(net239),
    .A2(\adder/adder/_0293_ ),
    .ZN(\adder/adder/_0014_ ));
 OAI21_X1 \adder/adder/_1931_  (.A(\adder/adder/_0014_ ),
    .B1(net214),
    .B2(net239),
    .ZN(\adder/adder/_0015_ ));
 XNOR2_X2 \adder/adder/_1932_  (.A(\adder/adder/_0864_ ),
    .B(\adder/adder/_0015_ ),
    .ZN(\adder/adder/_0016_ ));
 XNOR2_X2 \adder/adder/_1933_  (.A(\adder/adder/_0013_ ),
    .B(\adder/adder/_0016_ ),
    .ZN(\adder/adder/_0017_ ));
 NAND2_X1 \adder/adder/_1934_  (.A1(\adder/adder/_1037_ ),
    .A2(net252),
    .ZN(\adder/adder/_0018_ ));
 NAND2_X1 \adder/adder/_1935_  (.A1(\adder/adder/_1041_ ),
    .A2(\adder/adder/_0421_ ),
    .ZN(\adder/adder/_0019_ ));
 NAND3_X1 \adder/adder/_1936_  (.A1(\adder/adder/_0018_ ),
    .A2(\adder/adder/_0443_ ),
    .A3(\adder/adder/_0019_ ),
    .ZN(\adder/adder/_0020_ ));
 XNOR2_X2 \adder/adder/_1937_  (.A(\adder/adder/_0020_ ),
    .B(\adder/adder/_0766_ ),
    .ZN(\adder/adder/_0021_ ));
 NAND2_X1 \adder/adder/_1938_  (.A1(net239),
    .A2(\adder/adder/_0272_ ),
    .ZN(\adder/adder/_0022_ ));
 OAI21_X1 \adder/adder/_1939_  (.A(\adder/adder/_0022_ ),
    .B1(net215),
    .B2(net239),
    .ZN(\adder/adder/_0023_ ));
 XNOR2_X2 \adder/adder/_1940_  (.A(\adder/adder/_0864_ ),
    .B(\adder/adder/_0023_ ),
    .ZN(\adder/adder/_0024_ ));
 XNOR2_X2 \adder/adder/_1941_  (.A(\adder/adder/_0021_ ),
    .B(\adder/adder/_0024_ ),
    .ZN(\adder/adder/_0025_ ));
 NOR2_X1 \adder/adder/_1942_  (.A1(\adder/adder/_0017_ ),
    .A2(\adder/adder/_0025_ ),
    .ZN(\adder/adder/_0026_ ));
 NAND2_X1 \adder/adder/_1943_  (.A1(\adder/adder/_0967_ ),
    .A2(net252),
    .ZN(\adder/adder/_0027_ ));
 NAND2_X1 \adder/adder/_1944_  (.A1(\adder/adder/_0974_ ),
    .A2(\adder/adder/_0421_ ),
    .ZN(\adder/adder/_0028_ ));
 NAND3_X1 \adder/adder/_1945_  (.A1(\adder/adder/_0027_ ),
    .A2(\adder/adder/_0443_ ),
    .A3(\adder/adder/_0028_ ),
    .ZN(\adder/adder/_0029_ ));
 XNOR2_X2 \adder/adder/_1946_  (.A(\adder/adder/_0029_ ),
    .B(\adder/adder/_0766_ ),
    .ZN(\adder/adder/_0030_ ));
 NAND2_X1 \adder/adder/_1947_  (.A1(net239),
    .A2(\adder/adder/_0266_ ),
    .ZN(\adder/adder/_0031_ ));
 OAI21_X1 \adder/adder/_1948_  (.A(\adder/adder/_0031_ ),
    .B1(net216),
    .B2(net239),
    .ZN(\adder/adder/_0032_ ));
 XNOR2_X2 \adder/adder/_1949_  (.A(\adder/adder/_0864_ ),
    .B(\adder/adder/_0032_ ),
    .ZN(\adder/adder/_0033_ ));
 XNOR2_X2 \adder/adder/_1950_  (.A(\adder/adder/_0030_ ),
    .B(\adder/adder/_0033_ ),
    .ZN(\adder/adder/_0034_ ));
 NAND2_X1 \adder/adder/_1951_  (.A1(\adder/adder/_0986_ ),
    .A2(net252),
    .ZN(\adder/adder/_0035_ ));
 NAND2_X1 \adder/adder/_1952_  (.A1(\adder/adder/_0989_ ),
    .A2(\adder/adder/_0421_ ),
    .ZN(\adder/adder/_0036_ ));
 NAND3_X1 \adder/adder/_1953_  (.A1(\adder/adder/_0035_ ),
    .A2(\adder/adder/_0443_ ),
    .A3(\adder/adder/_0036_ ),
    .ZN(\adder/adder/_0037_ ));
 XNOR2_X1 \adder/adder/_1954_  (.A(\adder/adder/_0037_ ),
    .B(\adder/adder/_0766_ ),
    .ZN(\adder/adder/_0038_ ));
 NAND2_X1 \adder/adder/_1955_  (.A1(net239),
    .A2(net20),
    .ZN(\adder/adder/_0039_ ));
 OAI21_X1 \adder/adder/_1956_  (.A(\adder/adder/_0039_ ),
    .B1(\adder/adder/_0261_ ),
    .B2(net239),
    .ZN(\adder/adder/_0040_ ));
 XNOR2_X2 \adder/adder/_1957_  (.A(\adder/adder/_0863_ ),
    .B(\adder/adder/_0040_ ),
    .ZN(\adder/adder/_0041_ ));
 XNOR2_X1 \adder/adder/_1958_  (.A(\adder/adder/_0038_ ),
    .B(\adder/adder/_0041_ ),
    .ZN(\adder/adder/_0042_ ));
 NOR2_X1 \adder/adder/_1959_  (.A1(\adder/adder/_0034_ ),
    .A2(\adder/adder/_0042_ ),
    .ZN(\adder/adder/_0043_ ));
 NAND2_X1 \adder/adder/_1960_  (.A1(\adder/adder/_0026_ ),
    .A2(\adder/adder/_0043_ ),
    .ZN(\adder/adder/_0044_ ));
 NOR2_X1 \adder/adder/_1961_  (.A1(\adder/adder/_0009_ ),
    .A2(\adder/adder/_0044_ ),
    .ZN(\adder/adder/_0045_ ));
 NAND2_X1 \adder/adder/_1962_  (.A1(\adder/adder/_1063_ ),
    .A2(\adder/adder/_0045_ ),
    .ZN(\adder/adder/_0046_ ));
 NOR2_X1 \adder/adder/_1963_  (.A1(\adder/adder/_0021_ ),
    .A2(\adder/adder/_0024_ ),
    .ZN(\adder/adder/_0047_ ));
 INV_X1 \adder/adder/_1964_  (.A(\adder/adder/_0047_ ),
    .ZN(\adder/adder/_0048_ ));
 OR2_X1 \adder/adder/_1965_  (.A1(\adder/adder/_0013_ ),
    .A2(\adder/adder/_0016_ ),
    .ZN(\adder/adder/_0049_ ));
 OAI21_X1 \adder/adder/_1966_  (.A(\adder/adder/_0048_ ),
    .B1(\adder/adder/_0049_ ),
    .B2(\adder/adder/_0025_ ),
    .ZN(\adder/adder/_0051_ ));
 NAND2_X1 \adder/adder/_1967_  (.A1(\adder/adder/_0051_ ),
    .A2(\adder/adder/_0043_ ),
    .ZN(\adder/adder/_0052_ ));
 NOR2_X1 \adder/adder/_1968_  (.A1(\adder/adder/_0038_ ),
    .A2(\adder/adder/_0041_ ),
    .ZN(\adder/adder/_0053_ ));
 INV_X1 \adder/adder/_1969_  (.A(\adder/adder/_0042_ ),
    .ZN(\adder/adder/_0054_ ));
 NOR2_X1 \adder/adder/_1970_  (.A1(\adder/adder/_0030_ ),
    .A2(\adder/adder/_0033_ ),
    .ZN(\adder/adder/_0055_ ));
 AOI21_X1 \adder/adder/_1971_  (.A(\adder/adder/_0053_ ),
    .B1(\adder/adder/_0054_ ),
    .B2(\adder/adder/_0055_ ),
    .ZN(\adder/adder/_0056_ ));
 NAND2_X1 \adder/adder/_1972_  (.A1(\adder/adder/_0052_ ),
    .A2(\adder/adder/_0056_ ),
    .ZN(\adder/adder/_0057_ ));
 INV_X1 \adder/adder/_1973_  (.A(\adder/adder/_1092_ ),
    .ZN(\adder/adder/_0058_ ));
 OR2_X1 \adder/adder/_1974_  (.A1(\adder/adder/_1077_ ),
    .A2(\adder/adder/_1080_ ),
    .ZN(\adder/adder/_0059_ ));
 OAI21_X1 \adder/adder/_1975_  (.A(\adder/adder/_0058_ ),
    .B1(\adder/adder/_0059_ ),
    .B2(\adder/adder/_1091_ ),
    .ZN(\adder/adder/_0060_ ));
 NAND2_X1 \adder/adder/_1976_  (.A1(\adder/adder/_0060_ ),
    .A2(\adder/adder/_0008_ ),
    .ZN(\adder/adder/_0062_ ));
 OR2_X1 \adder/adder/_1977_  (.A1(\adder/adder/_1102_ ),
    .A2(\adder/adder/_1105_ ),
    .ZN(\adder/adder/_0063_ ));
 NOR2_X1 \adder/adder/_1978_  (.A1(\adder/adder/_0063_ ),
    .A2(\adder/adder/_0007_ ),
    .ZN(\adder/adder/_0064_ ));
 NOR2_X1 \adder/adder/_1979_  (.A1(\adder/adder/_0003_ ),
    .A2(\adder/adder/_0006_ ),
    .ZN(\adder/adder/_0065_ ));
 NOR2_X1 \adder/adder/_1980_  (.A1(\adder/adder/_0064_ ),
    .A2(\adder/adder/_0065_ ),
    .ZN(\adder/adder/_0066_ ));
 NAND2_X1 \adder/adder/_1981_  (.A1(\adder/adder/_0062_ ),
    .A2(\adder/adder/_0066_ ),
    .ZN(\adder/adder/_0067_ ));
 INV_X1 \adder/adder/_1982_  (.A(\adder/adder/_0044_ ),
    .ZN(\adder/adder/_0068_ ));
 AOI21_X1 \adder/adder/_1983_  (.A(\adder/adder/_0057_ ),
    .B1(\adder/adder/_0067_ ),
    .B2(\adder/adder/_0068_ ),
    .ZN(\adder/adder/_0069_ ));
 NAND2_X2 \adder/adder/_1984_  (.A1(\adder/adder/_0046_ ),
    .A2(\adder/adder/_0069_ ),
    .ZN(\adder/adder/_0070_ ));
 NAND2_X1 \adder/adder/_1985_  (.A1(net239),
    .A2(\adder/adder/_0322_ ),
    .ZN(\adder/adder/_0071_ ));
 OAI21_X1 \adder/adder/_1986_  (.A(\adder/adder/_0071_ ),
    .B1(\operand_fp16_fp32[19] ),
    .B2(net239),
    .ZN(\adder/adder/_0073_ ));
 XNOR2_X1 \adder/adder/_1987_  (.A(\adder/adder/_0864_ ),
    .B(\adder/adder/_0073_ ),
    .ZN(\adder/adder/_0074_ ));
 NAND3_X1 \adder/adder/_1988_  (.A1(\adder/adder/_0975_ ),
    .A2(net253),
    .A3(net252),
    .ZN(\adder/adder/_0075_ ));
 BUF_X1 input36 (.A(operand_fp32_i[27]),
    .Z(net36));
 XNOR2_X1 \adder/adder/_1990_  (.A(\adder/adder/_0075_ ),
    .B(\adder/adder/_0766_ ),
    .ZN(\adder/adder/_0077_ ));
 OR2_X1 \adder/adder/_1991_  (.A1(\adder/adder/_0074_ ),
    .A2(\adder/adder/_0077_ ),
    .ZN(\adder/adder/_0078_ ));
 NAND2_X1 \adder/adder/_1992_  (.A1(\adder/adder/_0074_ ),
    .A2(\adder/adder/_0077_ ),
    .ZN(\adder/adder/_0079_ ));
 NAND2_X2 \adder/adder/_1993_  (.A1(\adder/adder/_0078_ ),
    .A2(\adder/adder/_0079_ ),
    .ZN(\adder/adder/_0080_ ));
 BUF_X1 input35 (.A(operand_fp32_i[26]),
    .Z(net35));
 NAND3_X1 \adder/adder/_1995_  (.A1(\adder/adder/_0990_ ),
    .A2(net253),
    .A3(net252),
    .ZN(\adder/adder/_0082_ ));
 XNOR2_X2 \adder/adder/_1996_  (.A(\adder/adder/_0767_ ),
    .B(\adder/adder/_0082_ ),
    .ZN(\adder/adder/_0084_ ));
 NAND2_X1 \adder/adder/_1997_  (.A1(net239),
    .A2(\adder/adder/_0315_ ),
    .ZN(\adder/adder/_0085_ ));
 OAI21_X1 \adder/adder/_1998_  (.A(\adder/adder/_0085_ ),
    .B1(\operand_fp16_fp32[20] ),
    .B2(net239),
    .ZN(\adder/adder/_0086_ ));
 XNOR2_X2 \adder/adder/_1999_  (.A(\adder/adder/_0863_ ),
    .B(\adder/adder/_0086_ ),
    .ZN(\adder/adder/_0087_ ));
 XNOR2_X2 \adder/adder/_2000_  (.A(\adder/adder/_0084_ ),
    .B(\adder/adder/_0087_ ),
    .ZN(\adder/adder/_0088_ ));
 NOR2_X1 \adder/adder/_2001_  (.A1(\adder/adder/_0080_ ),
    .A2(\adder/adder/_0088_ ),
    .ZN(\adder/adder/_0089_ ));
 NAND3_X1 \adder/adder/_2002_  (.A1(\adder/adder/_1021_ ),
    .A2(net253),
    .A3(net252),
    .ZN(\adder/adder/_0090_ ));
 XNOR2_X2 \adder/adder/_2003_  (.A(\adder/adder/_0090_ ),
    .B(\adder/adder/_0766_ ),
    .ZN(\adder/adder/_0091_ ));
 NAND2_X1 \adder/adder/_2004_  (.A1(\adder/adder/_0414_ ),
    .A2(\adder/adder/_0319_ ),
    .ZN(\adder/adder/_0092_ ));
 OAI21_X1 \adder/adder/_2005_  (.A(\adder/adder/_0092_ ),
    .B1(net25),
    .B2(\adder/adder/_0414_ ),
    .ZN(\adder/adder/_0093_ ));
 XNOR2_X2 \adder/adder/_2006_  (.A(\adder/adder/_0864_ ),
    .B(\adder/adder/_0093_ ),
    .ZN(\adder/adder/_0095_ ));
 XNOR2_X2 \adder/adder/_2007_  (.A(\adder/adder/_0091_ ),
    .B(\adder/adder/_0095_ ),
    .ZN(\adder/adder/_0096_ ));
 NAND2_X1 \adder/adder/_2008_  (.A1(\adder/adder/_1043_ ),
    .A2(net253),
    .ZN(\adder/adder/_0097_ ));
 XNOR2_X1 \adder/adder/_2009_  (.A(\adder/adder/_0097_ ),
    .B(\adder/adder/_0766_ ),
    .ZN(\adder/adder/_0098_ ));
 NAND2_X1 \adder/adder/_2010_  (.A1(\adder/adder/_0414_ ),
    .A2(\operand_fp16_fp32[18] ),
    .ZN(\adder/adder/_0099_ ));
 OAI21_X1 \adder/adder/_2011_  (.A(\adder/adder/_0099_ ),
    .B1(\adder/adder/_0326_ ),
    .B2(\adder/adder/_0414_ ),
    .ZN(\adder/adder/_0100_ ));
 XNOR2_X1 \adder/adder/_2012_  (.A(\adder/adder/_0863_ ),
    .B(\adder/adder/_0100_ ),
    .ZN(\adder/adder/_0101_ ));
 XNOR2_X1 \adder/adder/_2013_  (.A(\adder/adder/_0098_ ),
    .B(\adder/adder/_0101_ ),
    .ZN(\adder/adder/_0102_ ));
 NOR2_X1 \adder/adder/_2014_  (.A1(\adder/adder/_0096_ ),
    .A2(\adder/adder/_0102_ ),
    .ZN(\adder/adder/_0103_ ));
 AND2_X1 \adder/adder/_2015_  (.A1(\adder/adder/_0089_ ),
    .A2(\adder/adder/_0103_ ),
    .ZN(\adder/adder/_0104_ ));
 NAND2_X1 \adder/adder/_2016_  (.A1(\adder/adder/_1069_ ),
    .A2(net252),
    .ZN(\adder/adder/_0106_ ));
 NAND2_X1 \adder/adder/_2017_  (.A1(\adder/adder/_1073_ ),
    .A2(\adder/adder/_0421_ ),
    .ZN(\adder/adder/_0107_ ));
 NAND3_X1 \adder/adder/_2018_  (.A1(\adder/adder/_0106_ ),
    .A2(net253),
    .A3(\adder/adder/_0107_ ),
    .ZN(\adder/adder/_0108_ ));
 XNOR2_X2 \adder/adder/_2019_  (.A(\adder/adder/_0108_ ),
    .B(\adder/adder/_0766_ ),
    .ZN(\adder/adder/_0109_ ));
 NAND2_X1 \adder/adder/_2020_  (.A1(net239),
    .A2(\adder/adder/_0284_ ),
    .ZN(\adder/adder/_0110_ ));
 OAI21_X1 \adder/adder/_2021_  (.A(\adder/adder/_0110_ ),
    .B1(\operand_fp16_fp32[13] ),
    .B2(net239),
    .ZN(\adder/adder/_0111_ ));
 XNOR2_X2 \adder/adder/_2022_  (.A(\adder/adder/_0864_ ),
    .B(\adder/adder/_0111_ ),
    .ZN(\adder/adder/_0112_ ));
 XNOR2_X2 \adder/adder/_2023_  (.A(\adder/adder/_0109_ ),
    .B(\adder/adder/_0112_ ),
    .ZN(\adder/adder/_0113_ ));
 NAND2_X1 \adder/adder/_2024_  (.A1(\adder/adder/_0859_ ),
    .A2(net253),
    .ZN(\adder/adder/_0114_ ));
 XNOR2_X1 \adder/adder/_2025_  (.A(\adder/adder/_0114_ ),
    .B(\adder/adder/_0766_ ),
    .ZN(\adder/adder/_0115_ ));
 NAND2_X1 \adder/adder/_2026_  (.A1(net239),
    .A2(\adder/adder/_0253_ ),
    .ZN(\adder/adder/_0117_ ));
 OAI21_X1 \adder/adder/_2027_  (.A(\adder/adder/_0117_ ),
    .B1(\operand_fp16_fp32[14] ),
    .B2(net239),
    .ZN(\adder/adder/_0118_ ));
 XNOR2_X1 \adder/adder/_2028_  (.A(\adder/adder/_0864_ ),
    .B(\adder/adder/_0118_ ),
    .ZN(\adder/adder/_0119_ ));
 XNOR2_X1 \adder/adder/_2029_  (.A(\adder/adder/_0115_ ),
    .B(\adder/adder/_0119_ ),
    .ZN(\adder/adder/_0120_ ));
 NOR2_X1 \adder/adder/_2030_  (.A1(\adder/adder/_0113_ ),
    .A2(\adder/adder/_0120_ ),
    .ZN(\adder/adder/_0121_ ));
 NAND2_X1 \adder/adder/_2031_  (.A1(\adder/adder/_0922_ ),
    .A2(net253),
    .ZN(\adder/adder/_0122_ ));
 XNOR2_X1 \adder/adder/_2032_  (.A(\adder/adder/_0122_ ),
    .B(\adder/adder/_0766_ ),
    .ZN(\adder/adder/_0123_ ));
 NAND2_X1 \adder/adder/_2033_  (.A1(net239),
    .A2(\adder/adder/_0251_ ),
    .ZN(\adder/adder/_0124_ ));
 OAI21_X1 \adder/adder/_2034_  (.A(\adder/adder/_0124_ ),
    .B1(\operand_fp16_fp32[15] ),
    .B2(net239),
    .ZN(\adder/adder/_0125_ ));
 XNOR2_X2 \adder/adder/_2035_  (.A(\adder/adder/_0864_ ),
    .B(\adder/adder/_0125_ ),
    .ZN(\adder/adder/_0126_ ));
 XNOR2_X2 \adder/adder/_2036_  (.A(\adder/adder/_0123_ ),
    .B(\adder/adder/_0126_ ),
    .ZN(\adder/adder/_0128_ ));
 NAND2_X1 \adder/adder/_2037_  (.A1(\adder/adder/_0949_ ),
    .A2(net253),
    .ZN(\adder/adder/_0129_ ));
 XNOR2_X1 \adder/adder/_2038_  (.A(\adder/adder/_0129_ ),
    .B(\adder/adder/_0766_ ),
    .ZN(\adder/adder/_0130_ ));
 NAND2_X1 \adder/adder/_2039_  (.A1(net239),
    .A2(\adder/adder/_0331_ ),
    .ZN(\adder/adder/_0131_ ));
 OAI21_X1 \adder/adder/_2040_  (.A(\adder/adder/_0131_ ),
    .B1(\operand_fp16_fp32[16] ),
    .B2(net239),
    .ZN(\adder/adder/_0132_ ));
 XNOR2_X2 \adder/adder/_2041_  (.A(\adder/adder/_0864_ ),
    .B(\adder/adder/_0132_ ),
    .ZN(\adder/adder/_0133_ ));
 XNOR2_X2 \adder/adder/_2042_  (.A(\adder/adder/_0130_ ),
    .B(\adder/adder/_0133_ ),
    .ZN(\adder/adder/_0134_ ));
 NOR2_X1 \adder/adder/_2043_  (.A1(\adder/adder/_0128_ ),
    .A2(\adder/adder/_0134_ ),
    .ZN(\adder/adder/_0135_ ));
 NAND2_X1 \adder/adder/_2044_  (.A1(\adder/adder/_0121_ ),
    .A2(\adder/adder/_0135_ ),
    .ZN(\adder/adder/_0136_ ));
 INV_X1 \adder/adder/_2045_  (.A(\adder/adder/_0136_ ),
    .ZN(\adder/adder/_0137_ ));
 NAND3_X1 \adder/adder/_2046_  (.A1(\adder/adder/_0070_ ),
    .A2(\adder/adder/_0104_ ),
    .A3(\adder/adder/_0137_ ),
    .ZN(\adder/adder/_0139_ ));
 NAND2_X1 \adder/adder/_2047_  (.A1(\adder/adder/_0084_ ),
    .A2(\adder/adder/_0087_ ),
    .ZN(\adder/adder/_0140_ ));
 NOR2_X1 \adder/adder/_2048_  (.A1(\adder/adder/_0098_ ),
    .A2(\adder/adder/_0101_ ),
    .ZN(\adder/adder/_0141_ ));
 INV_X1 \adder/adder/_2049_  (.A(\adder/adder/_0102_ ),
    .ZN(\adder/adder/_0142_ ));
 NOR2_X1 \adder/adder/_2050_  (.A1(\adder/adder/_0091_ ),
    .A2(\adder/adder/_0095_ ),
    .ZN(\adder/adder/_0143_ ));
 AOI21_X1 \adder/adder/_2051_  (.A(\adder/adder/_0141_ ),
    .B1(\adder/adder/_0142_ ),
    .B2(\adder/adder/_0143_ ),
    .ZN(\adder/adder/_0144_ ));
 INV_X1 \adder/adder/_2052_  (.A(\adder/adder/_0089_ ),
    .ZN(\adder/adder/_0145_ ));
 OAI221_X1 \adder/adder/_2053_  (.A(\adder/adder/_0140_ ),
    .B1(\adder/adder/_0088_ ),
    .B2(\adder/adder/_0078_ ),
    .C1(\adder/adder/_0144_ ),
    .C2(\adder/adder/_0145_ ),
    .ZN(\adder/adder/_0146_ ));
 OR2_X1 \adder/adder/_2054_  (.A1(\adder/adder/_0130_ ),
    .A2(\adder/adder/_0133_ ),
    .ZN(\adder/adder/_0147_ ));
 OR2_X1 \adder/adder/_2055_  (.A1(\adder/adder/_0123_ ),
    .A2(\adder/adder/_0126_ ),
    .ZN(\adder/adder/_0148_ ));
 NOR2_X1 \adder/adder/_2056_  (.A1(\adder/adder/_0115_ ),
    .A2(\adder/adder/_0119_ ),
    .ZN(\adder/adder/_0150_ ));
 INV_X1 \adder/adder/_2057_  (.A(\adder/adder/_0120_ ),
    .ZN(\adder/adder/_0151_ ));
 NOR2_X1 \adder/adder/_2058_  (.A1(\adder/adder/_0109_ ),
    .A2(\adder/adder/_0112_ ),
    .ZN(\adder/adder/_0152_ ));
 AOI21_X1 \adder/adder/_2059_  (.A(\adder/adder/_0150_ ),
    .B1(\adder/adder/_0151_ ),
    .B2(\adder/adder/_0152_ ),
    .ZN(\adder/adder/_0153_ ));
 INV_X1 \adder/adder/_2060_  (.A(\adder/adder/_0135_ ),
    .ZN(\adder/adder/_0154_ ));
 OAI221_X2 \adder/adder/_2061_  (.A(\adder/adder/_0147_ ),
    .B1(\adder/adder/_0134_ ),
    .B2(\adder/adder/_0148_ ),
    .C1(\adder/adder/_0153_ ),
    .C2(\adder/adder/_0154_ ),
    .ZN(\adder/adder/_0155_ ));
 AOI21_X1 \adder/adder/_2062_  (.A(\adder/adder/_0146_ ),
    .B1(\adder/adder/_0155_ ),
    .B2(\adder/adder/_0104_ ),
    .ZN(\adder/adder/_0156_ ));
 NAND2_X1 \adder/adder/_2063_  (.A1(\adder/adder/_0139_ ),
    .A2(\adder/adder/_0156_ ),
    .ZN(\adder/adder/_0157_ ));
 NAND2_X1 \adder/adder/_2064_  (.A1(net239),
    .A2(\adder/adder/_0307_ ),
    .ZN(\adder/adder/_0158_ ));
 OAI21_X1 \adder/adder/_2065_  (.A(\adder/adder/_0158_ ),
    .B1(\operand_fp16_fp32[21] ),
    .B2(net239),
    .ZN(\adder/adder/_0159_ ));
 XNOR2_X2 \adder/adder/_2066_  (.A(\adder/adder/_0864_ ),
    .B(\adder/adder/_0159_ ),
    .ZN(\adder/adder/_0161_ ));
 NAND2_X1 \adder/adder/_2067_  (.A1(\adder/adder/_1074_ ),
    .A2(net253),
    .ZN(\adder/adder/_0162_ ));
 XNOR2_X2 \adder/adder/_2068_  (.A(\adder/adder/_0766_ ),
    .B(\adder/adder/_0162_ ),
    .ZN(\adder/adder/_0163_ ));
 XNOR2_X2 \adder/adder/_2069_  (.A(\adder/adder/_0161_ ),
    .B(\adder/adder/_0163_ ),
    .ZN(\adder/adder/_0164_ ));
 NAND2_X1 \adder/adder/_2070_  (.A1(\adder/adder/_0414_ ),
    .A2(\operand_fp16_fp32[22] ),
    .ZN(\adder/adder/_0165_ ));
 OAI21_X1 \adder/adder/_2071_  (.A(\adder/adder/_0165_ ),
    .B1(\adder/adder/_0302_ ),
    .B2(\adder/adder/_0414_ ),
    .ZN(\adder/adder/_0166_ ));
 XNOR2_X1 \adder/adder/_2072_  (.A(\adder/adder/_0863_ ),
    .B(\adder/adder/_0166_ ),
    .ZN(\adder/adder/_0167_ ));
 NAND3_X1 \adder/adder/_2073_  (.A1(\adder/adder/_0833_ ),
    .A2(net253),
    .A3(net252),
    .ZN(\adder/adder/_0168_ ));
 XNOR2_X1 \adder/adder/_2074_  (.A(\adder/adder/_0766_ ),
    .B(\adder/adder/_0168_ ),
    .ZN(\adder/adder/_0169_ ));
 XNOR2_X1 \adder/adder/_2075_  (.A(\adder/adder/_0167_ ),
    .B(\adder/adder/_0169_ ),
    .ZN(\adder/adder/_0170_ ));
 NOR2_X1 \adder/adder/_2076_  (.A1(\adder/adder/_0164_ ),
    .A2(\adder/adder/_0170_ ),
    .ZN(\adder/adder/_0172_ ));
 NAND2_X1 \adder/adder/_2077_  (.A1(\adder/adder/_0157_ ),
    .A2(\adder/adder/_0172_ ),
    .ZN(\adder/adder/_0173_ ));
 NOR2_X1 \adder/adder/_2078_  (.A1(\adder/adder/_0167_ ),
    .A2(\adder/adder/_0169_ ),
    .ZN(\adder/adder/_0174_ ));
 INV_X1 \adder/adder/_2079_  (.A(\adder/adder/_0170_ ),
    .ZN(\adder/adder/_0175_ ));
 NOR2_X1 \adder/adder/_2080_  (.A1(\adder/adder/_0161_ ),
    .A2(\adder/adder/_0163_ ),
    .ZN(\adder/adder/_0176_ ));
 AOI21_X1 \adder/adder/_2081_  (.A(\adder/adder/_0174_ ),
    .B1(\adder/adder/_0175_ ),
    .B2(\adder/adder/_0176_ ),
    .ZN(\adder/adder/_0177_ ));
 NAND2_X1 \adder/adder/_2082_  (.A1(\adder/adder/_0173_ ),
    .A2(\adder/adder/_0177_ ),
    .ZN(\adder/adder/_0178_ ));
 NAND2_X1 \adder/adder/_2083_  (.A1(net239),
    .A2(\adder/adder/_0338_ ),
    .ZN(\adder/adder/_0179_ ));
 OAI21_X1 \adder/adder/_2084_  (.A(\adder/adder/_0179_ ),
    .B1(\adder/hb_a_d ),
    .B2(net239),
    .ZN(\adder/adder/_0180_ ));
 XNOR2_X1 \adder/adder/_2085_  (.A(\adder/adder/_0864_ ),
    .B(\adder/adder/_0180_ ),
    .ZN(\adder/adder/_0181_ ));
 NAND2_X1 \adder/adder/_2086_  (.A1(\adder/adder/_1099_ ),
    .A2(net253),
    .ZN(\adder/adder/_0183_ ));
 XNOR2_X2 \adder/adder/_2087_  (.A(\adder/adder/_0766_ ),
    .B(\adder/adder/_0183_ ),
    .ZN(\adder/adder/_0184_ ));
 XNOR2_X2 \adder/adder/_2088_  (.A(\adder/adder/_0181_ ),
    .B(\adder/adder/_0184_ ),
    .ZN(\adder/adder/_0185_ ));
 INV_X1 \adder/adder/_2089_  (.A(\adder/adder/_0185_ ),
    .ZN(\adder/adder/_0186_ ));
 NAND2_X1 \adder/adder/_2090_  (.A1(\adder/adder/_0178_ ),
    .A2(\adder/adder/_0186_ ),
    .ZN(\adder/adder/_0187_ ));
 OR2_X1 \adder/adder/_2091_  (.A1(\adder/adder/_0181_ ),
    .A2(\adder/adder/_0184_ ),
    .ZN(\adder/adder/_0188_ ));
 AOI21_X4 \adder/adder/_2092_  (.A(\adder/adder/_0495_ ),
    .B1(\adder/adder/_0187_ ),
    .B2(\adder/adder/_0188_ ),
    .ZN(\adder/mant_prenorm_d[47] ));
 AND2_X2 \adder/adder/_2093_  (.A1(\adder/adder/_0765_ ),
    .A2(\adder/adder/_0777_ ),
    .ZN(\adder/mant_prenorm_d[20] ));
 NAND2_X1 \adder/adder/_2094_  (.A1(\adder/adder/_0778_ ),
    .A2(\adder/adder/_0495_ ),
    .ZN(\adder/adder/_0189_ ));
 XNOR2_X2 \adder/adder/_2095_  (.A(\adder/adder/_0189_ ),
    .B(\adder/adder/_0867_ ),
    .ZN(\adder/mant_prenorm_d[21] ));
 NAND3_X1 \adder/adder/_2096_  (.A1(\adder/adder/_0778_ ),
    .A2(\adder/adder/_0495_ ),
    .A3(\adder/adder/_0867_ ),
    .ZN(\adder/adder/_0191_ ));
 XOR2_X2 \adder/adder/_2097_  (.A(\adder/adder/_0191_ ),
    .B(\adder/adder/_0927_ ),
    .Z(\adder/mant_prenorm_d[22] ));
 NOR2_X1 \adder/adder/_2098_  (.A1(\adder/adder/_0191_ ),
    .A2(\adder/adder/_0927_ ),
    .ZN(\adder/adder/_0192_ ));
 XNOR2_X2 \adder/adder/_2099_  (.A(\adder/adder/_0192_ ),
    .B(\adder/adder/_0962_ ),
    .ZN(\adder/mant_prenorm_d[23] ));
 XNOR2_X2 \adder/adder/_2100_  (.A(\adder/adder/_0965_ ),
    .B(\adder/adder/_1032_ ),
    .ZN(\adder/mant_prenorm_d[24] ));
 NAND3_X1 \adder/adder/_2101_  (.A1(\adder/adder/_0965_ ),
    .A2(\adder/adder/_1030_ ),
    .A3(\adder/adder/_1031_ ),
    .ZN(\adder/adder/_0193_ ));
 NAND2_X1 \adder/adder/_2102_  (.A1(\adder/adder/_0193_ ),
    .A2(\adder/adder/_1030_ ),
    .ZN(\adder/adder/_0194_ ));
 XNOR2_X2 \adder/adder/_2103_  (.A(\adder/adder/_0194_ ),
    .B(\adder/adder/_1050_ ),
    .ZN(\adder/mant_prenorm_d[25] ));
 OAI21_X1 \adder/adder/_2104_  (.A(\adder/adder/_1060_ ),
    .B1(\adder/adder/_0193_ ),
    .B2(\adder/adder/_1050_ ),
    .ZN(\adder/adder/_0195_ ));
 XNOR2_X2 \adder/adder/_2105_  (.A(\adder/adder/_0195_ ),
    .B(\adder/adder/_0982_ ),
    .ZN(\adder/mant_prenorm_d[26] ));
 INV_X1 \adder/adder/_2106_  (.A(\adder/adder/_0982_ ),
    .ZN(\adder/adder/_0197_ ));
 AOI21_X1 \adder/adder/_2107_  (.A(\adder/adder/_1054_ ),
    .B1(\adder/adder/_0195_ ),
    .B2(\adder/adder/_0197_ ),
    .ZN(\adder/adder/_0198_ ));
 XOR2_X2 \adder/adder/_2108_  (.A(\adder/adder/_0198_ ),
    .B(\adder/adder/_1000_ ),
    .Z(\adder/mant_prenorm_d[27] ));
 XNOR2_X2 \adder/adder/_2109_  (.A(\adder/adder/_1063_ ),
    .B(\adder/adder/_1081_ ),
    .ZN(\adder/mant_prenorm_d[28] ));
 INV_X1 \adder/adder/_2110_  (.A(\adder/adder/_1063_ ),
    .ZN(\adder/adder/_0199_ ));
 OAI21_X1 \adder/adder/_2111_  (.A(\adder/adder/_0059_ ),
    .B1(\adder/adder/_0199_ ),
    .B2(\adder/adder/_1081_ ),
    .ZN(\adder/adder/_0200_ ));
 XNOR2_X2 \adder/adder/_2112_  (.A(\adder/adder/_0200_ ),
    .B(\adder/adder/_1093_ ),
    .ZN(\adder/mant_prenorm_d[29] ));
 AND2_X1 \adder/adder/_2113_  (.A1(\adder/adder/_1063_ ),
    .A2(\adder/adder/_1094_ ),
    .ZN(\adder/adder/_0201_ ));
 NOR2_X1 \adder/adder/_2114_  (.A1(\adder/adder/_0201_ ),
    .A2(\adder/adder/_0060_ ),
    .ZN(\adder/adder/_0202_ ));
 XOR2_X2 \adder/adder/_2115_  (.A(\adder/adder/_0202_ ),
    .B(\adder/adder/_1106_ ),
    .Z(\adder/mant_prenorm_d[30] ));
 OAI21_X1 \adder/adder/_2116_  (.A(\adder/adder/_0063_ ),
    .B1(\adder/adder/_0202_ ),
    .B2(\adder/adder/_1106_ ),
    .ZN(\adder/adder/_0204_ ));
 XNOR2_X2 \adder/adder/_2117_  (.A(\adder/adder/_0204_ ),
    .B(\adder/adder/_0007_ ),
    .ZN(\adder/mant_prenorm_d[31] ));
 INV_X1 \adder/adder/_2118_  (.A(\adder/adder/_0067_ ),
    .ZN(\adder/adder/_0205_ ));
 OAI21_X2 \adder/adder/_2119_  (.A(\adder/adder/_0205_ ),
    .B1(\adder/adder/_0199_ ),
    .B2(\adder/adder/_0009_ ),
    .ZN(\adder/adder/_0206_ ));
 XNOR2_X2 \adder/adder/_2120_  (.A(\adder/adder/_0206_ ),
    .B(\adder/adder/_0017_ ),
    .ZN(\adder/mant_prenorm_d[32] ));
 INV_X1 \adder/adder/_2121_  (.A(\adder/adder/_0017_ ),
    .ZN(\adder/adder/_0207_ ));
 NAND2_X1 \adder/adder/_2122_  (.A1(\adder/adder/_0206_ ),
    .A2(\adder/adder/_0207_ ),
    .ZN(\adder/adder/_0208_ ));
 NAND2_X1 \adder/adder/_2123_  (.A1(\adder/adder/_0208_ ),
    .A2(\adder/adder/_0049_ ),
    .ZN(\adder/adder/_0209_ ));
 XNOR2_X2 \adder/adder/_2124_  (.A(\adder/adder/_0209_ ),
    .B(\adder/adder/_0025_ ),
    .ZN(\adder/mant_prenorm_d[33] ));
 NAND2_X1 \adder/adder/_2125_  (.A1(\adder/adder/_0206_ ),
    .A2(\adder/adder/_0026_ ),
    .ZN(\adder/adder/_0210_ ));
 INV_X1 \adder/adder/_2126_  (.A(\adder/adder/_0051_ ),
    .ZN(\adder/adder/_0212_ ));
 NAND2_X1 \adder/adder/_2127_  (.A1(\adder/adder/_0210_ ),
    .A2(\adder/adder/_0212_ ),
    .ZN(\adder/adder/_0213_ ));
 XNOR2_X2 \adder/adder/_2128_  (.A(\adder/adder/_0213_ ),
    .B(\adder/adder/_0034_ ),
    .ZN(\adder/mant_prenorm_d[34] ));
 INV_X1 \adder/adder/_2129_  (.A(\adder/adder/_0034_ ),
    .ZN(\adder/adder/_0214_ ));
 AOI21_X1 \adder/adder/_2130_  (.A(\adder/adder/_0055_ ),
    .B1(\adder/adder/_0213_ ),
    .B2(\adder/adder/_0214_ ),
    .ZN(\adder/adder/_0215_ ));
 XNOR2_X2 \adder/adder/_2131_  (.A(\adder/adder/_0215_ ),
    .B(\adder/adder/_0054_ ),
    .ZN(\adder/mant_prenorm_d[35] ));
 XNOR2_X2 \adder/adder/_2132_  (.A(\adder/adder/_0070_ ),
    .B(\adder/adder/_0113_ ),
    .ZN(\adder/mant_prenorm_d[36] ));
 INV_X1 \adder/adder/_2133_  (.A(\adder/adder/_0113_ ),
    .ZN(\adder/adder/_0216_ ));
 AOI21_X1 \adder/adder/_2134_  (.A(\adder/adder/_0152_ ),
    .B1(\adder/adder/_0070_ ),
    .B2(\adder/adder/_0216_ ),
    .ZN(\adder/adder/_0217_ ));
 XNOR2_X2 \adder/adder/_2135_  (.A(\adder/adder/_0217_ ),
    .B(\adder/adder/_0151_ ),
    .ZN(\adder/mant_prenorm_d[37] ));
 NAND2_X1 \adder/adder/_2136_  (.A1(\adder/adder/_0070_ ),
    .A2(\adder/adder/_0121_ ),
    .ZN(\adder/adder/_0219_ ));
 NAND2_X1 \adder/adder/_2137_  (.A1(\adder/adder/_0219_ ),
    .A2(\adder/adder/_0153_ ),
    .ZN(\adder/adder/_0220_ ));
 XNOR2_X2 \adder/adder/_2138_  (.A(\adder/adder/_0220_ ),
    .B(\adder/adder/_0128_ ),
    .ZN(\adder/mant_prenorm_d[38] ));
 INV_X1 \adder/adder/_2139_  (.A(\adder/adder/_0220_ ),
    .ZN(\adder/adder/_0221_ ));
 OAI21_X1 \adder/adder/_2140_  (.A(\adder/adder/_0148_ ),
    .B1(\adder/adder/_0221_ ),
    .B2(\adder/adder/_0128_ ),
    .ZN(\adder/adder/_0222_ ));
 XNOR2_X2 \adder/adder/_2141_  (.A(\adder/adder/_0222_ ),
    .B(\adder/adder/_0134_ ),
    .ZN(\adder/mant_prenorm_d[39] ));
 NAND2_X1 \adder/adder/_2142_  (.A1(\adder/adder/_0070_ ),
    .A2(\adder/adder/_0137_ ),
    .ZN(\adder/adder/_0223_ ));
 INV_X1 \adder/adder/_2143_  (.A(\adder/adder/_0155_ ),
    .ZN(\adder/adder/_0224_ ));
 NAND2_X1 \adder/adder/_2144_  (.A1(\adder/adder/_0223_ ),
    .A2(\adder/adder/_0224_ ),
    .ZN(\adder/adder/_0225_ ));
 XNOR2_X2 \adder/adder/_2145_  (.A(\adder/adder/_0225_ ),
    .B(\adder/adder/_0096_ ),
    .ZN(\adder/mant_prenorm_d[40] ));
 INV_X1 \adder/adder/_2146_  (.A(\adder/adder/_0096_ ),
    .ZN(\adder/adder/_0227_ ));
 AOI21_X1 \adder/adder/_2147_  (.A(\adder/adder/_0143_ ),
    .B1(\adder/adder/_0225_ ),
    .B2(\adder/adder/_0227_ ),
    .ZN(\adder/adder/_0228_ ));
 XNOR2_X2 \adder/adder/_2148_  (.A(\adder/adder/_0228_ ),
    .B(\adder/adder/_0142_ ),
    .ZN(\adder/mant_prenorm_d[41] ));
 NAND2_X1 \adder/adder/_2149_  (.A1(\adder/adder/_0225_ ),
    .A2(\adder/adder/_0103_ ),
    .ZN(\adder/adder/_0229_ ));
 NAND2_X1 \adder/adder/_2150_  (.A1(\adder/adder/_0229_ ),
    .A2(\adder/adder/_0144_ ),
    .ZN(\adder/adder/_0230_ ));
 XNOR2_X2 \adder/adder/_2151_  (.A(\adder/adder/_0230_ ),
    .B(\adder/adder/_0080_ ),
    .ZN(\adder/mant_prenorm_d[42] ));
 INV_X1 \adder/adder/_2152_  (.A(\adder/adder/_0080_ ),
    .ZN(\adder/adder/_0231_ ));
 NAND2_X1 \adder/adder/_2153_  (.A1(\adder/adder/_0230_ ),
    .A2(\adder/adder/_0231_ ),
    .ZN(\adder/adder/_0232_ ));
 NAND2_X1 \adder/adder/_2154_  (.A1(\adder/adder/_0232_ ),
    .A2(\adder/adder/_0078_ ),
    .ZN(\adder/adder/_0233_ ));
 NAND2_X1 \adder/adder/_2155_  (.A1(\adder/adder/_0233_ ),
    .A2(\adder/adder/_0088_ ),
    .ZN(\adder/adder/_0234_ ));
 INV_X1 \adder/adder/_2156_  (.A(\adder/adder/_0088_ ),
    .ZN(\adder/adder/_0236_ ));
 NAND3_X1 \adder/adder/_2157_  (.A1(\adder/adder/_0232_ ),
    .A2(\adder/adder/_0236_ ),
    .A3(\adder/adder/_0078_ ),
    .ZN(\adder/adder/_0237_ ));
 NAND2_X2 \adder/adder/_2158_  (.A1(\adder/adder/_0234_ ),
    .A2(\adder/adder/_0237_ ),
    .ZN(\adder/mant_prenorm_d[43] ));
 XNOR2_X2 \adder/adder/_2159_  (.A(\adder/adder/_0157_ ),
    .B(\adder/adder/_0164_ ),
    .ZN(\adder/mant_prenorm_d[44] ));
 INV_X1 \adder/adder/_2160_  (.A(\adder/adder/_0164_ ),
    .ZN(\adder/adder/_0238_ ));
 AOI21_X1 \adder/adder/_2161_  (.A(\adder/adder/_0176_ ),
    .B1(\adder/adder/_0157_ ),
    .B2(\adder/adder/_0238_ ),
    .ZN(\adder/adder/_0239_ ));
 XNOR2_X2 \adder/adder/_2162_  (.A(\adder/adder/_0239_ ),
    .B(\adder/adder/_0175_ ),
    .ZN(\adder/mant_prenorm_d[45] ));
 XNOR2_X2 \adder/adder/_2163_  (.A(\adder/adder/_0178_ ),
    .B(\adder/adder/_0185_ ),
    .ZN(\adder/mant_prenorm_d[46] ));
 INV_X1 \adder/adder/_2164_  (.A(net217),
    .ZN(\adder/adder/_0050_ ));
 NAND2_X1 \adder/adder/_2165_  (.A1(\adder/adder/_0050_ ),
    .A2(net46),
    .ZN(\adder/adder/_0061_ ));
 INV_X1 \adder/adder/_2166_  (.A(net45),
    .ZN(\adder/adder/_0072_ ));
 NOR2_X1 \adder/adder/_2167_  (.A1(\adder/adder/_0072_ ),
    .A2(net218),
    .ZN(\adder/adder/_0083_ ));
 INV_X1 \adder/adder/_2168_  (.A(net219),
    .ZN(\adder/adder/_0094_ ));
 NAND2_X1 \adder/adder/_2169_  (.A1(\adder/adder/_0094_ ),
    .A2(net42),
    .ZN(\adder/adder/_0105_ ));
 INV_X1 \adder/adder/_2170_  (.A(net39),
    .ZN(\adder/adder/_0116_ ));
 NOR2_X1 \adder/adder/_2171_  (.A1(\adder/adder/_0116_ ),
    .A2(net220),
    .ZN(\adder/adder/_0127_ ));
 INV_X1 \adder/adder/_2172_  (.A(net221),
    .ZN(\adder/adder/_0138_ ));
 INV_X1 \adder/adder/_2173_  (.A(net222),
    .ZN(\adder/adder/_0149_ ));
 OAI22_X1 \adder/adder/_2174_  (.A1(\adder/adder/_0138_ ),
    .A2(net28),
    .B1(\adder/adder/_0149_ ),
    .B2(net17),
    .ZN(\adder/adder/_0160_ ));
 INV_X1 \adder/adder/_2175_  (.A(net28),
    .ZN(\adder/adder/_0171_ ));
 OAI21_X1 \adder/adder/_2176_  (.A(\adder/adder/_0160_ ),
    .B1(net223),
    .B2(\adder/adder/_0171_ ),
    .ZN(\adder/adder/_0182_ ));
 NAND2_X1 \adder/adder/_2177_  (.A1(\adder/adder/_0116_ ),
    .A2(net224),
    .ZN(\adder/adder/_0190_ ));
 AOI21_X1 \adder/adder/_2178_  (.A(\adder/adder/_0127_ ),
    .B1(\adder/adder/_0182_ ),
    .B2(\adder/adder/_0190_ ),
    .ZN(\adder/adder/_0196_ ));
 NOR2_X1 \adder/adder/_2179_  (.A1(\adder/adder/_0094_ ),
    .A2(net42),
    .ZN(\adder/adder/_0203_ ));
 OAI21_X1 \adder/adder/_2180_  (.A(\adder/adder/_0105_ ),
    .B1(\adder/adder/_0196_ ),
    .B2(\adder/adder/_0203_ ),
    .ZN(\adder/adder/_0211_ ));
 INV_X1 \adder/adder/_2181_  (.A(net225),
    .ZN(\adder/adder/_0218_ ));
 OAI21_X1 \adder/adder/_2182_  (.A(\adder/adder/_0211_ ),
    .B1(net43),
    .B2(\adder/adder/_0218_ ),
    .ZN(\adder/adder/_0226_ ));
 INV_X1 \adder/adder/_2183_  (.A(net43),
    .ZN(\adder/adder/_0235_ ));
 OAI21_X1 \adder/adder/_2184_  (.A(\adder/adder/_0226_ ),
    .B1(\adder/adder/_0235_ ),
    .B2(net226),
    .ZN(\adder/adder/_0240_ ));
 INV_X1 \adder/adder/_2185_  (.A(net44),
    .ZN(\adder/adder/_0241_ ));
 NAND2_X1 \adder/adder/_2186_  (.A1(\adder/adder/_0241_ ),
    .A2(net227),
    .ZN(\adder/adder/_0242_ ));
 NAND2_X1 \adder/adder/_2187_  (.A1(\adder/adder/_0240_ ),
    .A2(\adder/adder/_0242_ ),
    .ZN(\adder/adder/_0243_ ));
 INV_X1 \adder/adder/_2188_  (.A(net228),
    .ZN(\adder/adder/_0244_ ));
 NAND2_X1 \adder/adder/_2189_  (.A1(\adder/adder/_0244_ ),
    .A2(net44),
    .ZN(\adder/adder/_0245_ ));
 NAND2_X1 \adder/adder/_2190_  (.A1(\adder/adder/_0243_ ),
    .A2(\adder/adder/_0245_ ),
    .ZN(\adder/adder/_0246_ ));
 NAND2_X1 \adder/adder/_2191_  (.A1(\adder/adder/_0072_ ),
    .A2(net229),
    .ZN(\adder/adder/_0247_ ));
 AOI21_X1 \adder/adder/_2192_  (.A(\adder/adder/_0083_ ),
    .B1(\adder/adder/_0246_ ),
    .B2(\adder/adder/_0247_ ),
    .ZN(\adder/adder/_0248_ ));
 NOR2_X1 \adder/adder/_2193_  (.A1(\adder/adder/_0050_ ),
    .A2(net46),
    .ZN(\adder/adder/_0249_ ));
 OAI21_X1 \adder/adder/_2194_  (.A(\adder/adder/_0061_ ),
    .B1(\adder/adder/_0248_ ),
    .B2(\adder/adder/_0249_ ),
    .ZN(\adder/adder/_0250_ ));
 INV_X1 \adder/adder/_2195_  (.A(net23),
    .ZN(\adder/adder/_0251_ ));
 NOR2_X1 \adder/adder/_2196_  (.A1(\adder/adder/_0251_ ),
    .A2(\operand_fp16_fp32[15] ),
    .ZN(\adder/adder/_0252_ ));
 INV_X1 \adder/adder/_2197_  (.A(net22),
    .ZN(\adder/adder/_0253_ ));
 AND2_X1 \adder/adder/_2198_  (.A1(\adder/adder/_0253_ ),
    .A2(\operand_fp16_fp32[14] ),
    .ZN(\adder/adder/_0254_ ));
 INV_X1 \adder/adder/_2199_  (.A(\operand_fp16_fp32[15] ),
    .ZN(\adder/adder/_0255_ ));
 NOR2_X1 \adder/adder/_2200_  (.A1(\adder/adder/_0255_ ),
    .A2(net23),
    .ZN(\adder/adder/_0256_ ));
 NOR2_X1 \adder/adder/_2201_  (.A1(\adder/adder/_0253_ ),
    .A2(\operand_fp16_fp32[14] ),
    .ZN(\adder/adder/_0257_ ));
 NOR4_X2 \adder/adder/_2202_  (.A1(\adder/adder/_0252_ ),
    .A2(\adder/adder/_0254_ ),
    .A3(\adder/adder/_0256_ ),
    .A4(\adder/adder/_0257_ ),
    .ZN(\adder/adder/_0258_ ));
 BUF_X1 input34 (.A(operand_fp32_i[25]),
    .Z(net34));
 XNOR2_X1 \adder/adder/_2204_  (.A(\operand_fp16_fp32[13] ),
    .B(net21),
    .ZN(\adder/adder/_0260_ ));
 INV_X1 \adder/adder/_2205_  (.A(net230),
    .ZN(\adder/adder/_0261_ ));
 CLKBUF_X2 input33 (.A(operand_fp32_i[24]),
    .Z(net33));
 NAND2_X1 \adder/adder/_2207_  (.A1(\adder/adder/_0261_ ),
    .A2(net20),
    .ZN(\adder/adder/_0263_ ));
 OR2_X1 \adder/adder/_2208_  (.A1(\adder/adder/_0261_ ),
    .A2(net20),
    .ZN(\adder/adder/_0264_ ));
 NAND4_X2 \adder/adder/_2209_  (.A1(\adder/adder/_0258_ ),
    .A2(\adder/adder/_0260_ ),
    .A3(\adder/adder/_0263_ ),
    .A4(\adder/adder/_0264_ ),
    .ZN(\adder/adder/_0265_ ));
 INV_X1 \adder/adder/_2210_  (.A(net19),
    .ZN(\adder/adder/_0266_ ));
 NOR2_X1 \adder/adder/_2211_  (.A1(\adder/adder/_0266_ ),
    .A2(net231),
    .ZN(\adder/adder/_0267_ ));
 NAND2_X1 \adder/adder/_2212_  (.A1(\adder/adder/_0266_ ),
    .A2(net232),
    .ZN(\adder/adder/_0268_ ));
 INV_X1 \adder/adder/_2213_  (.A(\adder/adder/_0268_ ),
    .ZN(\adder/adder/_0269_ ));
 INV_X1 \adder/adder/_2214_  (.A(net233),
    .ZN(\adder/adder/_0270_ ));
 NOR2_X1 \adder/adder/_2215_  (.A1(\adder/adder/_0270_ ),
    .A2(net18),
    .ZN(\adder/adder/_0271_ ));
 INV_X1 \adder/adder/_2216_  (.A(net18),
    .ZN(\adder/adder/_0272_ ));
 NOR2_X1 \adder/adder/_2217_  (.A1(\adder/adder/_0272_ ),
    .A2(net234),
    .ZN(\adder/adder/_0273_ ));
 NOR4_X1 \adder/adder/_2218_  (.A1(\adder/adder/_0267_ ),
    .A2(\adder/adder/_0269_ ),
    .A3(\adder/adder/_0271_ ),
    .A4(\adder/adder/_0273_ ),
    .ZN(\adder/adder/_0274_ ));
 XNOR2_X1 \adder/adder/_2219_  (.A(net235),
    .B(net48),
    .ZN(\adder/adder/_0275_ ));
 INV_X1 \adder/adder/_2220_  (.A(net236),
    .ZN(\adder/adder/_0276_ ));
 NAND2_X1 \adder/adder/_2221_  (.A1(\adder/adder/_0276_ ),
    .A2(net47),
    .ZN(\adder/adder/_0277_ ));
 INV_X1 \adder/adder/_2222_  (.A(net47),
    .ZN(\adder/adder/_0278_ ));
 NAND2_X1 \adder/adder/_2223_  (.A1(\adder/adder/_0278_ ),
    .A2(net237),
    .ZN(\adder/adder/_0279_ ));
 NAND4_X1 \adder/adder/_2224_  (.A1(\adder/adder/_0274_ ),
    .A2(\adder/adder/_0275_ ),
    .A3(\adder/adder/_0277_ ),
    .A4(\adder/adder/_0279_ ),
    .ZN(\adder/adder/_0280_ ));
 NOR2_X1 \adder/adder/_2225_  (.A1(\adder/adder/_0265_ ),
    .A2(\adder/adder/_0280_ ),
    .ZN(\adder/adder/_0281_ ));
 NAND2_X1 \adder/adder/_2226_  (.A1(\adder/adder/_0250_ ),
    .A2(\adder/adder/_0281_ ),
    .ZN(\adder/adder/_0282_ ));
 NAND3_X1 \adder/adder/_2227_  (.A1(\adder/adder/_0260_ ),
    .A2(net20),
    .A3(\adder/adder/_0261_ ),
    .ZN(\adder/adder/_0283_ ));
 INV_X1 \adder/adder/_2228_  (.A(net21),
    .ZN(\adder/adder/_0284_ ));
 OAI21_X1 \adder/adder/_2229_  (.A(\adder/adder/_0283_ ),
    .B1(\operand_fp16_fp32[13] ),
    .B2(\adder/adder/_0284_ ),
    .ZN(\adder/adder/_0285_ ));
 NAND2_X1 \adder/adder/_2230_  (.A1(\adder/adder/_0258_ ),
    .A2(\adder/adder/_0285_ ),
    .ZN(\adder/adder/_0286_ ));
 INV_X1 \adder/adder/_2231_  (.A(\adder/adder/_0256_ ),
    .ZN(\adder/adder/_0287_ ));
 AOI21_X1 \adder/adder/_2232_  (.A(\adder/adder/_0252_ ),
    .B1(\adder/adder/_0287_ ),
    .B2(\adder/adder/_0257_ ),
    .ZN(\adder/adder/_0288_ ));
 NAND2_X1 \adder/adder/_2233_  (.A1(\adder/adder/_0286_ ),
    .A2(\adder/adder/_0288_ ),
    .ZN(\adder/adder/_0289_ ));
 INV_X1 \adder/adder/_2234_  (.A(\adder/adder/_0289_ ),
    .ZN(\adder/adder/_0290_ ));
 INV_X1 \adder/adder/_2235_  (.A(\adder/adder/_0265_ ),
    .ZN(\adder/adder/_0291_ ));
 NAND3_X1 \adder/adder/_2236_  (.A1(\adder/adder/_0275_ ),
    .A2(net47),
    .A3(\adder/adder/_0276_ ),
    .ZN(\adder/adder/_0292_ ));
 INV_X1 \adder/adder/_2237_  (.A(net48),
    .ZN(\adder/adder/_0293_ ));
 OAI21_X1 \adder/adder/_2238_  (.A(\adder/adder/_0292_ ),
    .B1(net238),
    .B2(\adder/adder/_0293_ ),
    .ZN(\adder/adder/_0294_ ));
 NAND2_X1 \adder/adder/_2239_  (.A1(\adder/adder/_0274_ ),
    .A2(\adder/adder/_0294_ ),
    .ZN(\adder/adder/_0295_ ));
 AOI21_X1 \adder/adder/_2240_  (.A(\adder/adder/_0267_ ),
    .B1(\adder/adder/_0268_ ),
    .B2(\adder/adder/_0273_ ),
    .ZN(\adder/adder/_0296_ ));
 NAND2_X1 \adder/adder/_2241_  (.A1(\adder/adder/_0295_ ),
    .A2(\adder/adder/_0296_ ),
    .ZN(\adder/adder/_0297_ ));
 NAND2_X1 \adder/adder/_2242_  (.A1(\adder/adder/_0291_ ),
    .A2(\adder/adder/_0297_ ),
    .ZN(\adder/adder/_0298_ ));
 NAND3_X1 \adder/adder/_2243_  (.A1(\adder/adder/_0282_ ),
    .A2(\adder/adder/_0290_ ),
    .A3(\adder/adder/_0298_ ),
    .ZN(\adder/adder/_0299_ ));
 BUF_X1 input32 (.A(operand_fp32_i[23]),
    .Z(net32));
 XNOR2_X1 \adder/adder/_2245_  (.A(\adder/hb_b_d ),
    .B(\adder/hb_a_d ),
    .ZN(\adder/adder/_0301_ ));
 INV_X1 \adder/adder/_2246_  (.A(net31),
    .ZN(\adder/adder/_0302_ ));
 NOR2_X1 \adder/adder/_2247_  (.A1(\adder/adder/_0302_ ),
    .A2(\operand_fp16_fp32[22] ),
    .ZN(\adder/adder/_0303_ ));
 INV_X1 \adder/adder/_2248_  (.A(\adder/adder/_0303_ ),
    .ZN(\adder/adder/_0304_ ));
 NAND2_X1 \adder/adder/_2249_  (.A1(\adder/adder/_0302_ ),
    .A2(\operand_fp16_fp32[22] ),
    .ZN(\adder/adder/_0305_ ));
 NAND3_X1 \adder/adder/_2250_  (.A1(\adder/adder/_0301_ ),
    .A2(\adder/adder/_0304_ ),
    .A3(\adder/adder/_0305_ ),
    .ZN(\adder/adder/_0306_ ));
 INV_X1 \adder/adder/_2251_  (.A(net30),
    .ZN(\adder/adder/_0307_ ));
 LOGIC0_X1 \adder/adder/_1317__202  (.Z(net202));
 BUF_X1 input31 (.A(operand_fp32_i[22]),
    .Z(net31));
 BUF_X1 input30 (.A(operand_fp32_i[21]),
    .Z(net30));
 BUF_X1 input29 (.A(operand_fp32_i[20]),
    .Z(net29));
 BUF_X1 input28 (.A(operand_fp32_i[1]),
    .Z(net28));
 BUF_X1 input27 (.A(operand_fp32_i[19]),
    .Z(net27));
 BUF_X1 input26 (.A(operand_fp32_i[18]),
    .Z(net26));
 BUF_X1 input25 (.A(operand_fp32_i[17]),
    .Z(net25));
 BUF_X1 input24 (.A(operand_fp32_i[16]),
    .Z(net24));
 BUF_X1 input23 (.A(operand_fp32_i[15]),
    .Z(net23));
 BUF_X1 input22 (.A(operand_fp32_i[14]),
    .Z(net22));
 BUF_X1 input21 (.A(operand_fp32_i[13]),
    .Z(net21));
 BUF_X1 input20 (.A(operand_fp32_i[12]),
    .Z(net20));
 BUF_X1 input19 (.A(operand_fp32_i[11]),
    .Z(net19));
 BUF_X1 input18 (.A(operand_fp32_i[10]),
    .Z(net18));
 BUF_X1 input17 (.A(operand_fp32_i[0]),
    .Z(net17));
 BUF_X1 input16 (.A(operand_fp16_i[9]),
    .Z(net16));
 BUF_X1 input15 (.A(operand_fp16_i[8]),
    .Z(net15));
 BUF_X1 input14 (.A(operand_fp16_i[7]),
    .Z(net14));
 BUF_X1 input13 (.A(operand_fp16_i[6]),
    .Z(net13));
 BUF_X1 input12 (.A(operand_fp16_i[5]),
    .Z(net12));
 BUF_X2 input11 (.A(operand_fp16_i[4]),
    .Z(net11));
 BUF_X1 input10 (.A(operand_fp16_i[3]),
    .Z(net10));
 NOR2_X1 \adder/norm/LOD/_157_  (.A1(\adder/mant_prenorm_d[46] ),
    .A2(\adder/mant_prenorm_d[47] ),
    .ZN(\adder/norm/LOD/_113_ ));
 NOR2_X1 \adder/norm/LOD/_158_  (.A1(\adder/mant_prenorm_d[44] ),
    .A2(\adder/mant_prenorm_d[45] ),
    .ZN(\adder/norm/LOD/_114_ ));
 NAND2_X2 \adder/norm/LOD/_159_  (.A1(\adder/norm/LOD/_113_ ),
    .A2(\adder/norm/LOD/_114_ ),
    .ZN(\adder/norm/LOD/_115_ ));
 INV_X1 \adder/norm/LOD/_160_  (.A(\adder/norm/LOD/_115_ ),
    .ZN(\adder/norm/LOD/_116_ ));
 INV_X1 \adder/norm/LOD/_161_  (.A(\adder/mant_prenorm_d[42] ),
    .ZN(\adder/norm/LOD/_117_ ));
 AOI21_X1 \adder/norm/LOD/_162_  (.A(\adder/mant_prenorm_d[43] ),
    .B1(\adder/norm/LOD/_117_ ),
    .B2(\adder/mant_prenorm_d[41] ),
    .ZN(\adder/norm/LOD/_118_ ));
 NAND2_X1 \adder/norm/LOD/_163_  (.A1(\adder/norm/LOD/_116_ ),
    .A2(\adder/norm/LOD/_118_ ),
    .ZN(\adder/norm/LOD/_119_ ));
 INV_X1 \adder/norm/LOD/_164_  (.A(\adder/mant_prenorm_d[46] ),
    .ZN(\adder/norm/LOD/_120_ ));
 AOI21_X1 \adder/norm/LOD/_165_  (.A(\adder/mant_prenorm_d[47] ),
    .B1(\adder/norm/LOD/_120_ ),
    .B2(\adder/mant_prenorm_d[45] ),
    .ZN(\adder/norm/LOD/_121_ ));
 NAND2_X1 \adder/norm/LOD/_166_  (.A1(\adder/norm/LOD/_115_ ),
    .A2(\adder/norm/LOD/_121_ ),
    .ZN(\adder/norm/LOD/_122_ ));
 NAND2_X1 \adder/norm/LOD/_167_  (.A1(\adder/norm/LOD/_119_ ),
    .A2(\adder/norm/LOD/_122_ ),
    .ZN(\adder/norm/LOD/_123_ ));
 NOR2_X1 \adder/norm/LOD/_168_  (.A1(\adder/mant_prenorm_d[40] ),
    .A2(\adder/mant_prenorm_d[41] ),
    .ZN(\adder/norm/LOD/_124_ ));
 NOR2_X2 \adder/norm/LOD/_169_  (.A1(\adder/mant_prenorm_d[42] ),
    .A2(\adder/mant_prenorm_d[43] ),
    .ZN(\adder/norm/LOD/_125_ ));
 NAND2_X2 \adder/norm/LOD/_170_  (.A1(\adder/norm/LOD/_124_ ),
    .A2(\adder/norm/LOD/_125_ ),
    .ZN(\adder/norm/LOD/_126_ ));
 NOR2_X4 \adder/norm/LOD/_171_  (.A1(\adder/norm/LOD/_115_ ),
    .A2(\adder/norm/LOD/_126_ ),
    .ZN(\adder/norm/LOD/_127_ ));
 INV_X1 \adder/norm/LOD/_172_  (.A(\adder/norm/LOD/_127_ ),
    .ZN(\adder/norm/LOD/_128_ ));
 NAND2_X1 \adder/norm/LOD/_173_  (.A1(\adder/norm/LOD/_123_ ),
    .A2(\adder/norm/LOD/_128_ ),
    .ZN(\adder/norm/LOD/_129_ ));
 NOR2_X1 \adder/norm/LOD/_174_  (.A1(\adder/mant_prenorm_d[38] ),
    .A2(\adder/mant_prenorm_d[39] ),
    .ZN(\adder/norm/LOD/_130_ ));
 NOR2_X1 \adder/norm/LOD/_175_  (.A1(\adder/mant_prenorm_d[36] ),
    .A2(\adder/mant_prenorm_d[37] ),
    .ZN(\adder/norm/LOD/_131_ ));
 NAND2_X1 \adder/norm/LOD/_176_  (.A1(\adder/norm/LOD/_130_ ),
    .A2(\adder/norm/LOD/_131_ ),
    .ZN(\adder/norm/LOD/_132_ ));
 INV_X1 \adder/norm/LOD/_177_  (.A(\adder/norm/LOD/_132_ ),
    .ZN(\adder/norm/LOD/_133_ ));
 INV_X1 \adder/norm/LOD/_178_  (.A(\adder/mant_prenorm_d[34] ),
    .ZN(\adder/norm/LOD/_134_ ));
 AOI21_X1 \adder/norm/LOD/_179_  (.A(\adder/mant_prenorm_d[35] ),
    .B1(\adder/norm/LOD/_134_ ),
    .B2(\adder/mant_prenorm_d[33] ),
    .ZN(\adder/norm/LOD/_135_ ));
 NAND2_X1 \adder/norm/LOD/_180_  (.A1(\adder/norm/LOD/_133_ ),
    .A2(\adder/norm/LOD/_135_ ),
    .ZN(\adder/norm/LOD/_136_ ));
 INV_X1 \adder/norm/LOD/_181_  (.A(\adder/mant_prenorm_d[38] ),
    .ZN(\adder/norm/LOD/_137_ ));
 AOI21_X1 \adder/norm/LOD/_182_  (.A(\adder/mant_prenorm_d[39] ),
    .B1(\adder/norm/LOD/_137_ ),
    .B2(\adder/mant_prenorm_d[37] ),
    .ZN(\adder/norm/LOD/_138_ ));
 NAND2_X1 \adder/norm/LOD/_183_  (.A1(\adder/norm/LOD/_132_ ),
    .A2(\adder/norm/LOD/_138_ ),
    .ZN(\adder/norm/LOD/_139_ ));
 NAND2_X1 \adder/norm/LOD/_184_  (.A1(\adder/norm/LOD/_136_ ),
    .A2(\adder/norm/LOD/_139_ ),
    .ZN(\adder/norm/LOD/_140_ ));
 NAND2_X1 \adder/norm/LOD/_185_  (.A1(\adder/norm/LOD/_140_ ),
    .A2(\adder/norm/LOD/_127_ ),
    .ZN(\adder/norm/LOD/_141_ ));
 NAND2_X1 \adder/norm/LOD/_186_  (.A1(\adder/norm/LOD/_129_ ),
    .A2(\adder/norm/LOD/_141_ ),
    .ZN(\adder/norm/LOD/_142_ ));
 NOR2_X1 \adder/norm/LOD/_187_  (.A1(\adder/mant_prenorm_d[32] ),
    .A2(\adder/mant_prenorm_d[33] ),
    .ZN(\adder/norm/LOD/_143_ ));
 NOR2_X1 \adder/norm/LOD/_188_  (.A1(\adder/mant_prenorm_d[34] ),
    .A2(\adder/mant_prenorm_d[35] ),
    .ZN(\adder/norm/LOD/_144_ ));
 NAND2_X1 \adder/norm/LOD/_189_  (.A1(\adder/norm/LOD/_143_ ),
    .A2(\adder/norm/LOD/_144_ ),
    .ZN(\adder/norm/LOD/_145_ ));
 NOR2_X2 \adder/norm/LOD/_190_  (.A1(\adder/norm/LOD/_132_ ),
    .A2(\adder/norm/LOD/_145_ ),
    .ZN(\adder/norm/LOD/_146_ ));
 NAND2_X4 \adder/norm/LOD/_191_  (.A1(\adder/norm/LOD/_127_ ),
    .A2(\adder/norm/LOD/_146_ ),
    .ZN(\adder/norm/LOD/_147_ ));
 NAND2_X1 \adder/norm/LOD/_192_  (.A1(\adder/norm/LOD/_142_ ),
    .A2(\adder/norm/LOD/_147_ ),
    .ZN(\adder/norm/LOD/_148_ ));
 NOR2_X1 \adder/norm/LOD/_193_  (.A1(\adder/mant_prenorm_d[30] ),
    .A2(\adder/mant_prenorm_d[31] ),
    .ZN(\adder/norm/LOD/_149_ ));
 NOR2_X1 \adder/norm/LOD/_194_  (.A1(\adder/mant_prenorm_d[28] ),
    .A2(\adder/mant_prenorm_d[29] ),
    .ZN(\adder/norm/LOD/_150_ ));
 NAND2_X1 \adder/norm/LOD/_195_  (.A1(\adder/norm/LOD/_149_ ),
    .A2(\adder/norm/LOD/_150_ ),
    .ZN(\adder/norm/LOD/_151_ ));
 INV_X1 \adder/norm/LOD/_196_  (.A(\adder/norm/LOD/_151_ ),
    .ZN(\adder/norm/LOD/_152_ ));
 INV_X1 \adder/norm/LOD/_197_  (.A(\adder/mant_prenorm_d[26] ),
    .ZN(\adder/norm/LOD/_153_ ));
 AOI21_X1 \adder/norm/LOD/_198_  (.A(\adder/mant_prenorm_d[27] ),
    .B1(\adder/norm/LOD/_153_ ),
    .B2(\adder/mant_prenorm_d[25] ),
    .ZN(\adder/norm/LOD/_154_ ));
 NAND2_X1 \adder/norm/LOD/_199_  (.A1(\adder/norm/LOD/_152_ ),
    .A2(\adder/norm/LOD/_154_ ),
    .ZN(\adder/norm/LOD/_155_ ));
 INV_X1 \adder/norm/LOD/_200_  (.A(\adder/mant_prenorm_d[30] ),
    .ZN(\adder/norm/LOD/_156_ ));
 AOI21_X1 \adder/norm/LOD/_201_  (.A(\adder/mant_prenorm_d[31] ),
    .B1(\adder/norm/LOD/_156_ ),
    .B2(\adder/mant_prenorm_d[29] ),
    .ZN(\adder/norm/LOD/_000_ ));
 NAND2_X1 \adder/norm/LOD/_202_  (.A1(\adder/norm/LOD/_151_ ),
    .A2(\adder/norm/LOD/_000_ ),
    .ZN(\adder/norm/LOD/_001_ ));
 NAND2_X1 \adder/norm/LOD/_203_  (.A1(\adder/norm/LOD/_155_ ),
    .A2(\adder/norm/LOD/_001_ ),
    .ZN(\adder/norm/LOD/_002_ ));
 NOR2_X1 \adder/norm/LOD/_204_  (.A1(\adder/mant_prenorm_d[24] ),
    .A2(\adder/mant_prenorm_d[25] ),
    .ZN(\adder/norm/LOD/_003_ ));
 NOR2_X1 \adder/norm/LOD/_205_  (.A1(\adder/mant_prenorm_d[26] ),
    .A2(\adder/mant_prenorm_d[27] ),
    .ZN(\adder/norm/LOD/_004_ ));
 NAND2_X1 \adder/norm/LOD/_206_  (.A1(\adder/norm/LOD/_003_ ),
    .A2(\adder/norm/LOD/_004_ ),
    .ZN(\adder/norm/LOD/_005_ ));
 NOR2_X2 \adder/norm/LOD/_207_  (.A1(\adder/norm/LOD/_151_ ),
    .A2(\adder/norm/LOD/_005_ ),
    .ZN(\adder/norm/LOD/_006_ ));
 INV_X2 \adder/norm/LOD/_208_  (.A(\adder/norm/LOD/_006_ ),
    .ZN(\adder/norm/LOD/_007_ ));
 NAND2_X1 \adder/norm/LOD/_209_  (.A1(\adder/norm/LOD/_002_ ),
    .A2(\adder/norm/LOD/_007_ ),
    .ZN(\adder/norm/LOD/_008_ ));
 INV_X1 \adder/norm/LOD/_210_  (.A(\adder/mant_prenorm_d[22] ),
    .ZN(\adder/norm/LOD/_009_ ));
 INV_X1 \adder/norm/LOD/_211_  (.A(\adder/mant_prenorm_d[23] ),
    .ZN(\adder/norm/LOD/_010_ ));
 NAND2_X1 \adder/norm/LOD/_212_  (.A1(\adder/norm/LOD/_009_ ),
    .A2(\adder/norm/LOD/_010_ ),
    .ZN(\adder/norm/LOD/_011_ ));
 INV_X1 \adder/norm/LOD/_213_  (.A(\adder/mant_prenorm_d[20] ),
    .ZN(\adder/norm/LOD/_012_ ));
 INV_X1 \adder/norm/LOD/_214_  (.A(\adder/mant_prenorm_d[21] ),
    .ZN(\adder/norm/LOD/_013_ ));
 NAND2_X1 \adder/norm/LOD/_215_  (.A1(\adder/norm/LOD/_012_ ),
    .A2(\adder/norm/LOD/_013_ ),
    .ZN(\adder/norm/LOD/_014_ ));
 NOR2_X1 \adder/norm/LOD/_216_  (.A1(\adder/norm/LOD/_011_ ),
    .A2(\adder/norm/LOD/_014_ ),
    .ZN(\adder/norm/LOD/_015_ ));
 INV_X1 \adder/norm/LOD/_217_  (.A(net86),
    .ZN(\adder/norm/LOD/_016_ ));
 AOI21_X1 \adder/norm/LOD/_218_  (.A(net87),
    .B1(\adder/norm/LOD/_016_ ),
    .B2(net88),
    .ZN(\adder/norm/LOD/_017_ ));
 NAND2_X1 \adder/norm/LOD/_219_  (.A1(\adder/norm/LOD/_015_ ),
    .A2(\adder/norm/LOD/_017_ ),
    .ZN(\adder/norm/LOD/_018_ ));
 NOR2_X1 \adder/norm/LOD/_220_  (.A1(\adder/mant_prenorm_d[22] ),
    .A2(\adder/mant_prenorm_d[23] ),
    .ZN(\adder/norm/LOD/_019_ ));
 NOR2_X1 \adder/norm/LOD/_221_  (.A1(\adder/mant_prenorm_d[20] ),
    .A2(\adder/mant_prenorm_d[21] ),
    .ZN(\adder/norm/LOD/_020_ ));
 NAND2_X1 \adder/norm/LOD/_222_  (.A1(\adder/norm/LOD/_019_ ),
    .A2(\adder/norm/LOD/_020_ ),
    .ZN(\adder/norm/LOD/_021_ ));
 AOI21_X1 \adder/norm/LOD/_223_  (.A(\adder/mant_prenorm_d[23] ),
    .B1(\adder/norm/LOD/_009_ ),
    .B2(\adder/mant_prenorm_d[21] ),
    .ZN(\adder/norm/LOD/_022_ ));
 NAND2_X1 \adder/norm/LOD/_224_  (.A1(\adder/norm/LOD/_021_ ),
    .A2(\adder/norm/LOD/_022_ ),
    .ZN(\adder/norm/LOD/_023_ ));
 NAND2_X1 \adder/norm/LOD/_225_  (.A1(\adder/norm/LOD/_018_ ),
    .A2(\adder/norm/LOD/_023_ ),
    .ZN(\adder/norm/LOD/_024_ ));
 NAND2_X1 \adder/norm/LOD/_226_  (.A1(\adder/norm/LOD/_024_ ),
    .A2(\adder/norm/LOD/_006_ ),
    .ZN(\adder/norm/LOD/_025_ ));
 NAND2_X1 \adder/norm/LOD/_227_  (.A1(\adder/norm/LOD/_008_ ),
    .A2(\adder/norm/LOD/_025_ ),
    .ZN(\adder/norm/LOD/_026_ ));
 OR2_X2 \adder/norm/LOD/_228_  (.A1(net89),
    .A2(net90),
    .ZN(\adder/norm/LOD/_027_ ));
 INV_X1 \adder/norm/LOD/_229_  (.A(net91),
    .ZN(\adder/norm/LOD/_028_ ));
 INV_X1 \adder/norm/LOD/_230_  (.A(net92),
    .ZN(\adder/norm/LOD/_029_ ));
 NAND2_X1 \adder/norm/LOD/_231_  (.A1(\adder/norm/LOD/_028_ ),
    .A2(\adder/norm/LOD/_029_ ),
    .ZN(\adder/norm/LOD/_030_ ));
 NOR2_X1 \adder/norm/LOD/_232_  (.A1(\adder/norm/LOD/_027_ ),
    .A2(\adder/norm/LOD/_030_ ),
    .ZN(\adder/norm/LOD/_031_ ));
 NAND2_X1 \adder/norm/LOD/_233_  (.A1(\adder/norm/LOD/_031_ ),
    .A2(\adder/norm/LOD/_015_ ),
    .ZN(\adder/norm/LOD/_032_ ));
 NOR2_X1 \adder/norm/LOD/_234_  (.A1(\adder/norm/LOD/_007_ ),
    .A2(\adder/norm/LOD/_032_ ),
    .ZN(\adder/norm/LOD/_033_ ));
 NOR2_X2 \adder/norm/LOD/_235_  (.A1(\adder/norm/LOD/_033_ ),
    .A2(\adder/norm/LOD/_147_ ),
    .ZN(\adder/norm/Mant_leadingOne_D[4] ));
 NAND2_X1 \adder/norm/LOD/_236_  (.A1(\adder/norm/LOD/_026_ ),
    .A2(\adder/norm/Mant_leadingOne_D[4] ),
    .ZN(\adder/norm/LOD/_034_ ));
 NAND2_X1 \adder/norm/LOD/_237_  (.A1(\adder/norm/LOD/_148_ ),
    .A2(\adder/norm/LOD/_034_ ),
    .ZN(\adder/norm/LOD/_035_ ));
 INV_X1 \adder/norm/LOD/_238_  (.A(\adder/norm/LOD/_035_ ),
    .ZN(\adder/norm/LOD/_036_ ));
 NOR2_X2 \adder/norm/LOD/_239_  (.A1(net93),
    .A2(net94),
    .ZN(\adder/norm/LOD/_037_ ));
 INV_X1 \adder/norm/LOD/_240_  (.A(net95),
    .ZN(\adder/norm/LOD/_038_ ));
 INV_X1 \adder/norm/LOD/_241_  (.A(net96),
    .ZN(\adder/norm/LOD/_039_ ));
 NAND3_X2 \adder/norm/LOD/_242_  (.A1(\adder/norm/LOD/_037_ ),
    .A2(\adder/norm/LOD/_038_ ),
    .A3(\adder/norm/LOD/_039_ ),
    .ZN(\adder/norm/LOD/_040_ ));
 AOI21_X1 \adder/norm/LOD/_243_  (.A(net97),
    .B1(\adder/norm/LOD/_038_ ),
    .B2(net98),
    .ZN(\adder/norm/LOD/_041_ ));
 NAND2_X1 \adder/norm/LOD/_244_  (.A1(\adder/norm/LOD/_040_ ),
    .A2(\adder/norm/LOD/_041_ ),
    .ZN(\adder/norm/LOD/_042_ ));
 INV_X1 \adder/norm/LOD/_245_  (.A(net99),
    .ZN(\adder/norm/LOD/_043_ ));
 INV_X1 \adder/norm/LOD/_246_  (.A(net100),
    .ZN(\adder/norm/LOD/_044_ ));
 OAI21_X1 \adder/norm/LOD/_247_  (.A(\adder/norm/LOD/_043_ ),
    .B1(\adder/norm/LOD/_044_ ),
    .B2(net101),
    .ZN(\adder/norm/LOD/_045_ ));
 OAI21_X1 \adder/norm/LOD/_248_  (.A(\adder/norm/LOD/_042_ ),
    .B1(\adder/norm/LOD/_040_ ),
    .B2(\adder/norm/LOD/_045_ ),
    .ZN(\adder/norm/LOD/_046_ ));
 NOR2_X1 \adder/norm/LOD/_249_  (.A1(net102),
    .A2(net103),
    .ZN(\adder/norm/LOD/_047_ ));
 INV_X1 \adder/norm/LOD/_250_  (.A(net104),
    .ZN(\adder/norm/LOD/_048_ ));
 NAND3_X1 \adder/norm/LOD/_251_  (.A1(\adder/norm/LOD/_047_ ),
    .A2(\adder/norm/LOD/_048_ ),
    .A3(\adder/norm/LOD/_044_ ),
    .ZN(\adder/norm/LOD/_049_ ));
 NOR2_X2 \adder/norm/LOD/_252_  (.A1(\adder/norm/LOD/_049_ ),
    .A2(\adder/norm/LOD/_040_ ),
    .ZN(\adder/norm/LOD/_050_ ));
 INV_X1 \adder/norm/LOD/_253_  (.A(\adder/norm/LOD/_050_ ),
    .ZN(\adder/norm/LOD/_051_ ));
 NAND2_X1 \adder/norm/LOD/_254_  (.A1(\adder/norm/LOD/_046_ ),
    .A2(\adder/norm/LOD/_051_ ),
    .ZN(\adder/norm/LOD/_052_ ));
 NOR2_X2 \adder/norm/LOD/_255_  (.A1(net105),
    .A2(net106),
    .ZN(\adder/norm/LOD/_053_ ));
 INV_X1 \adder/norm/LOD/_256_  (.A(net107),
    .ZN(\adder/norm/LOD/_054_ ));
 INV_X1 \adder/norm/LOD/_257_  (.A(net108),
    .ZN(\adder/norm/LOD/_055_ ));
 NAND3_X1 \adder/norm/LOD/_258_  (.A1(\adder/norm/LOD/_053_ ),
    .A2(\adder/norm/LOD/_054_ ),
    .A3(\adder/norm/LOD/_055_ ),
    .ZN(\adder/norm/LOD/_056_ ));
 INV_X1 \adder/norm/LOD/_259_  (.A(net109),
    .ZN(\adder/norm/LOD/_057_ ));
 AOI21_X1 \adder/norm/LOD/_260_  (.A(net110),
    .B1(\adder/norm/LOD/_057_ ),
    .B2(net111),
    .ZN(\adder/norm/LOD/_058_ ));
 NAND2_X1 \adder/norm/LOD/_261_  (.A1(\adder/norm/LOD/_056_ ),
    .A2(\adder/norm/LOD/_058_ ),
    .ZN(\adder/norm/LOD/_059_ ));
 INV_X1 \adder/norm/LOD/_262_  (.A(net112),
    .ZN(\adder/norm/LOD/_060_ ));
 INV_X1 \adder/norm/LOD/_263_  (.A(net113),
    .ZN(\adder/norm/LOD/_061_ ));
 OAI21_X1 \adder/norm/LOD/_264_  (.A(\adder/norm/LOD/_060_ ),
    .B1(\adder/norm/LOD/_061_ ),
    .B2(net114),
    .ZN(\adder/norm/LOD/_062_ ));
 OAI21_X1 \adder/norm/LOD/_265_  (.A(\adder/norm/LOD/_059_ ),
    .B1(\adder/norm/LOD/_056_ ),
    .B2(\adder/norm/LOD/_062_ ),
    .ZN(\adder/norm/LOD/_063_ ));
 NAND2_X1 \adder/norm/LOD/_266_  (.A1(\adder/norm/LOD/_063_ ),
    .A2(\adder/norm/LOD/_050_ ),
    .ZN(\adder/norm/LOD/_064_ ));
 NAND2_X1 \adder/norm/LOD/_267_  (.A1(\adder/norm/LOD/_052_ ),
    .A2(\adder/norm/LOD/_064_ ),
    .ZN(\adder/norm/LOD/_065_ ));
 INV_X1 \adder/norm/LOD/_268_  (.A(\adder/norm/LOD/_056_ ),
    .ZN(\adder/norm/LOD/_066_ ));
 NOR2_X1 \adder/norm/LOD/_269_  (.A1(net115),
    .A2(net116),
    .ZN(\adder/norm/LOD/_067_ ));
 NOR2_X1 \adder/norm/LOD/_270_  (.A1(net117),
    .A2(net118),
    .ZN(\adder/norm/LOD/_068_ ));
 NAND3_X1 \adder/norm/LOD/_271_  (.A1(\adder/norm/LOD/_066_ ),
    .A2(\adder/norm/LOD/_067_ ),
    .A3(\adder/norm/LOD/_068_ ),
    .ZN(\adder/norm/LOD/_069_ ));
 NOR2_X2 \adder/norm/LOD/_272_  (.A1(\adder/norm/LOD/_069_ ),
    .A2(\adder/norm/LOD/_051_ ),
    .ZN(\adder/norm/LOD/_070_ ));
 INV_X4 \adder/norm/LOD/_273_  (.A(\adder/norm/LOD/_147_ ),
    .ZN(\adder/norm/LOD/_071_ ));
 NAND2_X2 \adder/norm/LOD/_274_  (.A1(\adder/norm/LOD/_033_ ),
    .A2(\adder/norm/LOD/_071_ ),
    .ZN(\adder/norm/LOD/_072_ ));
 NOR2_X4 \adder/norm/LOD/_275_  (.A1(\adder/norm/LOD/_070_ ),
    .A2(\adder/norm/LOD/_072_ ),
    .ZN(\adder/norm/Mant_leadingOne_D[5] ));
 NAND2_X1 \adder/norm/LOD/_276_  (.A1(\adder/norm/LOD/_065_ ),
    .A2(\adder/norm/Mant_leadingOne_D[5] ),
    .ZN(\adder/norm/LOD/_073_ ));
 NAND2_X2 \adder/norm/LOD/_277_  (.A1(\adder/norm/LOD/_036_ ),
    .A2(\adder/norm/LOD/_073_ ),
    .ZN(\adder/norm/Mant_leadingOne_D[0] ));
 INV_X1 \adder/norm/LOD/_278_  (.A(\adder/mant_prenorm_d[31] ),
    .ZN(\adder/norm/LOD/_074_ ));
 NAND2_X1 \adder/norm/LOD/_279_  (.A1(\adder/norm/LOD/_156_ ),
    .A2(\adder/norm/LOD/_074_ ),
    .ZN(\adder/norm/LOD/_075_ ));
 INV_X1 \adder/norm/LOD/_280_  (.A(\adder/norm/LOD/_004_ ),
    .ZN(\adder/norm/LOD/_076_ ));
 AOI21_X1 \adder/norm/LOD/_281_  (.A(\adder/norm/LOD/_075_ ),
    .B1(\adder/norm/LOD/_076_ ),
    .B2(\adder/norm/LOD/_150_ ),
    .ZN(\adder/norm/LOD/_077_ ));
 NAND2_X1 \adder/norm/LOD/_282_  (.A1(\adder/norm/LOD/_007_ ),
    .A2(\adder/norm/LOD/_077_ ),
    .ZN(\adder/norm/LOD/_078_ ));
 AOI21_X1 \adder/norm/LOD/_283_  (.A(\adder/norm/LOD/_011_ ),
    .B1(\adder/norm/LOD/_027_ ),
    .B2(\adder/norm/LOD/_020_ ),
    .ZN(\adder/norm/LOD/_079_ ));
 NAND2_X1 \adder/norm/LOD/_284_  (.A1(\adder/norm/LOD/_079_ ),
    .A2(\adder/norm/LOD/_006_ ),
    .ZN(\adder/norm/LOD/_080_ ));
 NAND2_X1 \adder/norm/LOD/_285_  (.A1(\adder/norm/LOD/_078_ ),
    .A2(\adder/norm/LOD/_080_ ),
    .ZN(\adder/norm/LOD/_081_ ));
 NAND2_X1 \adder/norm/LOD/_286_  (.A1(\adder/norm/LOD/_081_ ),
    .A2(\adder/norm/LOD/_071_ ),
    .ZN(\adder/norm/LOD/_082_ ));
 INV_X1 \adder/norm/LOD/_287_  (.A(\adder/mant_prenorm_d[36] ),
    .ZN(\adder/norm/LOD/_083_ ));
 INV_X1 \adder/norm/LOD/_288_  (.A(\adder/mant_prenorm_d[37] ),
    .ZN(\adder/norm/LOD/_084_ ));
 NAND2_X1 \adder/norm/LOD/_289_  (.A1(\adder/norm/LOD/_083_ ),
    .A2(\adder/norm/LOD/_084_ ),
    .ZN(\adder/norm/LOD/_085_ ));
 OAI21_X1 \adder/norm/LOD/_290_  (.A(\adder/norm/LOD/_130_ ),
    .B1(\adder/norm/LOD/_085_ ),
    .B2(\adder/norm/LOD/_144_ ),
    .ZN(\adder/norm/LOD/_086_ ));
 NAND2_X1 \adder/norm/LOD/_291_  (.A1(\adder/norm/LOD/_127_ ),
    .A2(\adder/norm/LOD/_086_ ),
    .ZN(\adder/norm/LOD/_087_ ));
 NAND2_X1 \adder/norm/LOD/_292_  (.A1(\adder/norm/LOD/_116_ ),
    .A2(\adder/norm/LOD/_125_ ),
    .ZN(\adder/norm/LOD/_088_ ));
 NAND2_X1 \adder/norm/LOD/_293_  (.A1(\adder/norm/LOD/_115_ ),
    .A2(\adder/norm/LOD/_113_ ),
    .ZN(\adder/norm/LOD/_089_ ));
 NAND2_X1 \adder/norm/LOD/_294_  (.A1(\adder/norm/LOD/_088_ ),
    .A2(\adder/norm/LOD/_089_ ),
    .ZN(\adder/norm/LOD/_090_ ));
 NAND3_X1 \adder/norm/LOD/_295_  (.A1(\adder/norm/LOD/_147_ ),
    .A2(\adder/norm/LOD/_087_ ),
    .A3(\adder/norm/LOD/_090_ ),
    .ZN(\adder/norm/LOD/_091_ ));
 NAND2_X1 \adder/norm/LOD/_296_  (.A1(\adder/norm/LOD/_082_ ),
    .A2(\adder/norm/LOD/_091_ ),
    .ZN(\adder/norm/LOD/_092_ ));
 NAND2_X1 \adder/norm/LOD/_297_  (.A1(\adder/norm/LOD/_092_ ),
    .A2(\adder/norm/LOD/_072_ ),
    .ZN(\adder/norm/LOD/_093_ ));
 NOR2_X1 \adder/norm/LOD/_298_  (.A1(\adder/norm/LOD/_040_ ),
    .A2(\adder/norm/LOD/_047_ ),
    .ZN(\adder/norm/LOD/_094_ ));
 NOR3_X1 \adder/norm/LOD/_299_  (.A1(\adder/norm/LOD/_094_ ),
    .A2(net119),
    .A3(net120),
    .ZN(\adder/norm/LOD/_095_ ));
 OAI21_X1 \adder/norm/LOD/_300_  (.A(\adder/norm/LOD/_053_ ),
    .B1(\adder/norm/LOD/_056_ ),
    .B2(\adder/norm/LOD/_067_ ),
    .ZN(\adder/norm/LOD/_096_ ));
 NAND2_X1 \adder/norm/LOD/_301_  (.A1(\adder/norm/LOD/_096_ ),
    .A2(\adder/norm/LOD/_050_ ),
    .ZN(\adder/norm/LOD/_097_ ));
 NAND2_X1 \adder/norm/LOD/_302_  (.A1(\adder/norm/LOD/_095_ ),
    .A2(\adder/norm/LOD/_097_ ),
    .ZN(\adder/norm/LOD/_098_ ));
 INV_X1 \adder/norm/LOD/_303_  (.A(\adder/norm/LOD/_098_ ),
    .ZN(\adder/norm/LOD/_099_ ));
 NAND2_X1 \adder/norm/LOD/_304_  (.A1(\adder/norm/LOD/_099_ ),
    .A2(\adder/norm/Mant_leadingOne_D[5] ),
    .ZN(\adder/norm/LOD/_100_ ));
 NAND2_X2 \adder/norm/LOD/_305_  (.A1(\adder/norm/LOD/_093_ ),
    .A2(\adder/norm/LOD/_100_ ),
    .ZN(\adder/norm/Mant_leadingOne_D[1] ));
 INV_X1 \adder/norm/LOD/_306_  (.A(\adder/norm/LOD/_126_ ),
    .ZN(\adder/norm/LOD/_101_ ));
 AOI21_X1 \adder/norm/LOD/_307_  (.A(\adder/norm/LOD/_115_ ),
    .B1(\adder/norm/LOD/_101_ ),
    .B2(\adder/norm/LOD/_132_ ),
    .ZN(\adder/norm/LOD/_102_ ));
 NAND2_X1 \adder/norm/LOD/_308_  (.A1(\adder/norm/LOD/_147_ ),
    .A2(\adder/norm/LOD/_102_ ),
    .ZN(\adder/norm/LOD/_103_ ));
 OAI21_X1 \adder/norm/LOD/_309_  (.A(\adder/norm/LOD/_152_ ),
    .B1(\adder/norm/LOD/_015_ ),
    .B2(\adder/norm/LOD/_005_ ),
    .ZN(\adder/norm/LOD/_104_ ));
 OAI21_X1 \adder/norm/LOD/_310_  (.A(\adder/norm/LOD/_103_ ),
    .B1(\adder/norm/LOD/_147_ ),
    .B2(\adder/norm/LOD/_104_ ),
    .ZN(\adder/norm/LOD/_105_ ));
 NAND2_X1 \adder/norm/LOD/_311_  (.A1(\adder/norm/LOD/_105_ ),
    .A2(\adder/norm/LOD/_072_ ),
    .ZN(\adder/norm/LOD/_106_ ));
 AOI21_X1 \adder/norm/LOD/_312_  (.A(\adder/norm/LOD/_040_ ),
    .B1(\adder/norm/LOD/_050_ ),
    .B2(\adder/norm/LOD/_056_ ),
    .ZN(\adder/norm/LOD/_107_ ));
 NAND2_X1 \adder/norm/LOD/_313_  (.A1(\adder/norm/Mant_leadingOne_D[5] ),
    .A2(\adder/norm/LOD/_107_ ),
    .ZN(\adder/norm/LOD/_108_ ));
 NAND2_X1 \adder/norm/LOD/_314_  (.A1(\adder/norm/LOD/_106_ ),
    .A2(\adder/norm/LOD/_108_ ),
    .ZN(\adder/norm/Mant_leadingOne_D[2] ));
 INV_X1 \adder/norm/LOD/_315_  (.A(\adder/norm/LOD/_146_ ),
    .ZN(\adder/norm/LOD/_109_ ));
 OAI21_X1 \adder/norm/LOD/_316_  (.A(\adder/norm/LOD/_127_ ),
    .B1(\adder/norm/LOD/_109_ ),
    .B2(\adder/norm/LOD/_006_ ),
    .ZN(\adder/norm/LOD/_110_ ));
 INV_X1 \adder/norm/LOD/_317_  (.A(\adder/norm/LOD/_072_ ),
    .ZN(\adder/norm/LOD/_111_ ));
 NAND2_X1 \adder/norm/LOD/_318_  (.A1(\adder/norm/LOD/_069_ ),
    .A2(\adder/norm/LOD/_050_ ),
    .ZN(\adder/norm/LOD/_112_ ));
 AOI21_X1 \adder/norm/LOD/_319_  (.A(\adder/norm/LOD/_110_ ),
    .B1(\adder/norm/LOD/_111_ ),
    .B2(\adder/norm/LOD/_112_ ),
    .ZN(\adder/norm/Mant_leadingOne_D[3] ));
 AND2_X1 \adder/norm/LOD/_320_  (.A1(\adder/norm/LOD/_111_ ),
    .A2(\adder/norm/LOD/_070_ ),
    .ZN(\adder/norm/Mant_zero_S ));
 INV_X1 \adder/norm/_1476_  (.A(\adder/exp_prenorm_d[1] ),
    .ZN(\adder/norm/_1464_ ));
 NAND2_X1 \adder/norm/_1477_  (.A1(\adder/norm/_1464_ ),
    .A2(\adder/norm/Mant_leadingOne_D[1] ),
    .ZN(\adder/norm/_1475_ ));
 NOR2_X1 \adder/norm/_1478_  (.A1(\adder/norm/_1464_ ),
    .A2(\adder/norm/Mant_leadingOne_D[1] ),
    .ZN(\adder/norm/_0010_ ));
 INV_X1 \adder/norm/_1479_  (.A(\adder/exp_prenorm_d[0] ),
    .ZN(\adder/norm/_0021_ ));
 BUF_X1 input9 (.A(operand_fp16_i[2]),
    .Z(net9));
 NOR2_X1 \adder/norm/_1481_  (.A1(\adder/norm/_0021_ ),
    .A2(\adder/norm/Mant_leadingOne_D[0] ),
    .ZN(\adder/norm/_0042_ ));
 OAI21_X1 \adder/norm/_1482_  (.A(\adder/norm/_1475_ ),
    .B1(\adder/norm/_0010_ ),
    .B2(\adder/norm/_0042_ ),
    .ZN(\adder/norm/_0051_ ));
 INV_X1 \adder/norm/_1483_  (.A(\adder/exp_prenorm_d[2] ),
    .ZN(\adder/norm/_0061_ ));
 NAND2_X1 \adder/norm/_1484_  (.A1(\adder/norm/_0061_ ),
    .A2(\adder/norm/Mant_leadingOne_D[2] ),
    .ZN(\adder/norm/_0071_ ));
 INV_X1 \adder/norm/_1485_  (.A(\adder/norm/Mant_leadingOne_D[2] ),
    .ZN(\adder/norm/_0080_ ));
 NAND2_X1 \adder/norm/_1486_  (.A1(\adder/norm/_0080_ ),
    .A2(\adder/exp_prenorm_d[2] ),
    .ZN(\adder/norm/_0090_ ));
 NAND2_X1 \adder/norm/_1487_  (.A1(\adder/norm/_0071_ ),
    .A2(\adder/norm/_0090_ ),
    .ZN(\adder/norm/_0101_ ));
 INV_X1 \adder/norm/_1488_  (.A(\adder/exp_prenorm_d[3] ),
    .ZN(\adder/norm/_0112_ ));
 NAND2_X1 \adder/norm/_1489_  (.A1(\adder/norm/_0112_ ),
    .A2(\adder/norm/Mant_leadingOne_D[3] ),
    .ZN(\adder/norm/_0123_ ));
 INV_X2 \adder/norm/_1490_  (.A(\adder/norm/Mant_leadingOne_D[3] ),
    .ZN(\adder/norm/_0134_ ));
 NAND2_X2 \adder/norm/_1491_  (.A1(\adder/norm/_0134_ ),
    .A2(\adder/exp_prenorm_d[3] ),
    .ZN(\adder/norm/_0145_ ));
 NAND2_X2 \adder/norm/_1492_  (.A1(\adder/norm/_0123_ ),
    .A2(\adder/norm/_0145_ ),
    .ZN(\adder/norm/_0156_ ));
 NOR2_X1 \adder/norm/_1493_  (.A1(\adder/norm/_0101_ ),
    .A2(\adder/norm/_0156_ ),
    .ZN(\adder/norm/_0167_ ));
 NAND2_X1 \adder/norm/_1494_  (.A1(\adder/norm/_0051_ ),
    .A2(\adder/norm/_0167_ ),
    .ZN(\adder/norm/_0178_ ));
 NOR2_X1 \adder/norm/_1495_  (.A1(\adder/norm/_0156_ ),
    .A2(\adder/norm/_0071_ ),
    .ZN(\adder/norm/_0189_ ));
 INV_X1 \adder/norm/_1496_  (.A(\adder/norm/_0123_ ),
    .ZN(\adder/norm/_0200_ ));
 NOR2_X1 \adder/norm/_1497_  (.A1(\adder/norm/_0189_ ),
    .A2(\adder/norm/_0200_ ),
    .ZN(\adder/norm/_0211_ ));
 NAND2_X1 \adder/norm/_1498_  (.A1(\adder/norm/_0178_ ),
    .A2(\adder/norm/_0211_ ),
    .ZN(\adder/norm/_0222_ ));
 INV_X1 \adder/norm/_1499_  (.A(\adder/exp_prenorm_d[7] ),
    .ZN(\adder/norm/_0233_ ));
 BUF_X1 input8 (.A(operand_fp16_i[1]),
    .Z(net8));
 XNOR2_X1 \adder/norm/_1501_  (.A(\adder/norm/_0233_ ),
    .B(\adder/norm/Mant_leadingOne_D[5] ),
    .ZN(\adder/norm/_0255_ ));
 BUF_X1 input7 (.A(operand_fp16_i[15]),
    .Z(net7));
 INV_X1 \adder/norm/_1503_  (.A(\adder/exp_prenorm_d[6] ),
    .ZN(\adder/norm/_0277_ ));
 NAND2_X1 \adder/norm/_1504_  (.A1(\adder/norm/_0277_ ),
    .A2(\adder/norm/Mant_leadingOne_D[5] ),
    .ZN(\adder/norm/_0288_ ));
 INV_X2 \adder/norm/_1505_  (.A(\adder/norm/Mant_leadingOne_D[5] ),
    .ZN(\adder/norm/_0299_ ));
 NAND2_X1 \adder/norm/_1506_  (.A1(\adder/norm/_0299_ ),
    .A2(\adder/exp_prenorm_d[6] ),
    .ZN(\adder/norm/_0310_ ));
 NAND2_X1 \adder/norm/_1507_  (.A1(\adder/norm/_0288_ ),
    .A2(\adder/norm/_0310_ ),
    .ZN(\adder/norm/_0321_ ));
 NOR2_X1 \adder/norm/_1508_  (.A1(\adder/norm/_0255_ ),
    .A2(\adder/norm/_0321_ ),
    .ZN(\adder/norm/_0332_ ));
 INV_X1 \adder/norm/_1509_  (.A(\adder/norm/_0332_ ),
    .ZN(\adder/norm/_0343_ ));
 INV_X1 \adder/norm/_1510_  (.A(\adder/exp_prenorm_d[4] ),
    .ZN(\adder/norm/_0354_ ));
 NAND2_X1 \adder/norm/_1511_  (.A1(\adder/norm/_0354_ ),
    .A2(\adder/norm/Mant_leadingOne_D[4] ),
    .ZN(\adder/norm/_0365_ ));
 INV_X1 \adder/norm/_1512_  (.A(\adder/norm/Mant_leadingOne_D[4] ),
    .ZN(\adder/norm/_0376_ ));
 NAND2_X1 \adder/norm/_1513_  (.A1(\adder/norm/_0376_ ),
    .A2(\adder/exp_prenorm_d[4] ),
    .ZN(\adder/norm/_0387_ ));
 AND2_X1 \adder/norm/_1514_  (.A1(\adder/norm/_0365_ ),
    .A2(\adder/norm/_0387_ ),
    .ZN(\adder/norm/_0398_ ));
 CLKBUF_X3 input6 (.A(operand_fp16_i[14]),
    .Z(net6));
 XNOR2_X1 \adder/norm/_1516_  (.A(\adder/exp_prenorm_d[5] ),
    .B(\adder/norm/Mant_leadingOne_D[5] ),
    .ZN(\adder/norm/_0420_ ));
 NAND2_X1 \adder/norm/_1517_  (.A1(\adder/norm/_0398_ ),
    .A2(\adder/norm/_0420_ ),
    .ZN(\adder/norm/_0431_ ));
 NOR2_X1 \adder/norm/_1518_  (.A1(\adder/norm/_0343_ ),
    .A2(\adder/norm/_0431_ ),
    .ZN(\adder/norm/_0442_ ));
 NAND2_X1 \adder/norm/_1519_  (.A1(\adder/norm/_0222_ ),
    .A2(\adder/norm/_0442_ ),
    .ZN(\adder/norm/_0453_ ));
 NAND2_X1 \adder/norm/_1520_  (.A1(\adder/exp_prenorm_d[7] ),
    .A2(\adder/exp_prenorm_d[6] ),
    .ZN(\adder/norm/_0464_ ));
 NAND2_X1 \adder/norm/_1521_  (.A1(\adder/norm/_0464_ ),
    .A2(\adder/norm/Mant_leadingOne_D[5] ),
    .ZN(\adder/norm/_0475_ ));
 INV_X1 \adder/norm/_1522_  (.A(\adder/norm/_0475_ ),
    .ZN(\adder/norm/_0486_ ));
 INV_X1 \adder/norm/_1523_  (.A(\adder/exp_prenorm_d[5] ),
    .ZN(\adder/norm/_0497_ ));
 NAND2_X1 \adder/norm/_1524_  (.A1(\adder/norm/_0497_ ),
    .A2(\adder/norm/Mant_leadingOne_D[5] ),
    .ZN(\adder/norm/_0508_ ));
 NOR2_X1 \adder/norm/_1525_  (.A1(\adder/norm/_0497_ ),
    .A2(\adder/norm/Mant_leadingOne_D[5] ),
    .ZN(\adder/norm/_0519_ ));
 OAI21_X1 \adder/norm/_1526_  (.A(\adder/norm/_0508_ ),
    .B1(\adder/norm/_0519_ ),
    .B2(\adder/norm/_0365_ ),
    .ZN(\adder/norm/_0530_ ));
 AOI21_X1 \adder/norm/_1527_  (.A(\adder/norm/_0486_ ),
    .B1(\adder/norm/_0332_ ),
    .B2(\adder/norm/_0530_ ),
    .ZN(\adder/norm/_0541_ ));
 NAND2_X1 \adder/norm/_1528_  (.A1(\adder/norm/_0453_ ),
    .A2(\adder/norm/_0541_ ),
    .ZN(\adder/norm/_0552_ ));
 NOR2_X1 \adder/norm/_1529_  (.A1(net121),
    .A2(\adder/norm/Mant_leadingOne_D[5] ),
    .ZN(\adder/norm/_0563_ ));
 NAND2_X1 \adder/norm/_1530_  (.A1(\adder/norm/_0552_ ),
    .A2(\adder/norm/_0563_ ),
    .ZN(\adder/norm/_0574_ ));
 INV_X1 \adder/norm/_1531_  (.A(net122),
    .ZN(\adder/norm/_0585_ ));
 NAND2_X1 \adder/norm/_1532_  (.A1(\adder/norm/_0574_ ),
    .A2(\adder/norm/_0585_ ),
    .ZN(\adder/norm/_0596_ ));
 NAND4_X1 \adder/norm/_1533_  (.A1(\adder/norm/_0453_ ),
    .A2(net123),
    .A3(\adder/norm/Mant_leadingOne_D[5] ),
    .A4(\adder/norm/_0541_ ),
    .ZN(\adder/norm/_0602_ ));
 NAND2_X4 \adder/norm/_1534_  (.A1(\adder/norm/_0596_ ),
    .A2(\adder/norm/_0602_ ),
    .ZN(\adder/norm/_0609_ ));
 INV_X2 \adder/norm/_1535_  (.A(\adder/norm/Mant_zero_S ),
    .ZN(\adder/norm/_0616_ ));
 NAND2_X4 \adder/norm/_1536_  (.A1(\adder/norm/_0616_ ),
    .A2(\adder/norm/_0609_ ),
    .ZN(\adder/norm/_0622_ ));
 NAND2_X1 \adder/norm/_1537_  (.A1(\adder/norm/_0622_ ),
    .A2(\adder/norm/_0354_ ),
    .ZN(\adder/norm/_0628_ ));
 NAND3_X1 \adder/norm/_1538_  (.A1(\adder/norm/_0609_ ),
    .A2(\adder/norm/_0376_ ),
    .A3(\adder/norm/_0616_ ),
    .ZN(\adder/norm/_0634_ ));
 NAND2_X1 \adder/norm/_1539_  (.A1(\adder/norm/_0628_ ),
    .A2(\adder/norm/_0634_ ),
    .ZN(\adder/norm/_0635_ ));
 NAND2_X1 \adder/norm/_1540_  (.A1(\adder/norm/_0622_ ),
    .A2(\adder/norm/_0061_ ),
    .ZN(\adder/norm/_0636_ ));
 NAND3_X1 \adder/norm/_1541_  (.A1(\adder/norm/_0609_ ),
    .A2(\adder/norm/_0080_ ),
    .A3(\adder/norm/_0616_ ),
    .ZN(\adder/norm/_0637_ ));
 NAND2_X4 \adder/norm/_1542_  (.A1(\adder/norm/_0637_ ),
    .A2(\adder/norm/_0636_ ),
    .ZN(\adder/norm/_0638_ ));
 BUF_X1 input5 (.A(operand_fp16_i[13]),
    .Z(net5));
 NAND2_X2 \adder/norm/_1544_  (.A1(\adder/norm/_0622_ ),
    .A2(\adder/norm/_0112_ ),
    .ZN(\adder/norm/_0640_ ));
 NAND3_X4 \adder/norm/_1545_  (.A1(\adder/norm/_0609_ ),
    .A2(\adder/norm/_0134_ ),
    .A3(\adder/norm/_0616_ ),
    .ZN(\adder/norm/_0641_ ));
 NAND2_X4 \adder/norm/_1546_  (.A1(\adder/norm/_0640_ ),
    .A2(\adder/norm/_0641_ ),
    .ZN(\adder/norm/_0642_ ));
 NAND3_X4 \adder/norm/_1547_  (.A1(\adder/norm/_0635_ ),
    .A2(\adder/norm/_0638_ ),
    .A3(\adder/norm/_0642_ ),
    .ZN(\adder/norm/_0643_ ));
 NAND2_X1 \adder/norm/_1548_  (.A1(net257),
    .A2(\adder/exp_prenorm_d[5] ),
    .ZN(\adder/norm/_0644_ ));
 OAI21_X4 \adder/norm/_1549_  (.A(\adder/norm/_0644_ ),
    .B1(\adder/norm/_0299_ ),
    .B2(net257),
    .ZN(\adder/norm/_0645_ ));
 INV_X4 \adder/norm/_1550_  (.A(\adder/norm/_0622_ ),
    .ZN(\adder/norm/_0646_ ));
 INV_X1 \adder/norm/_1551_  (.A(net124),
    .ZN(\adder/norm/_0647_ ));
 NOR2_X1 \adder/norm/_1552_  (.A1(\adder/norm/_0646_ ),
    .A2(\adder/norm/_0647_ ),
    .ZN(\adder/norm/_0648_ ));
 NOR2_X1 \adder/norm/_1553_  (.A1(\adder/norm/_0646_ ),
    .A2(\adder/norm/_0277_ ),
    .ZN(\adder/norm/_0649_ ));
 NOR2_X2 \adder/norm/_1554_  (.A1(\adder/norm/_0646_ ),
    .A2(\adder/norm/_0233_ ),
    .ZN(\adder/norm/_0650_ ));
 NAND2_X1 \adder/norm/_1555_  (.A1(\adder/norm/_0649_ ),
    .A2(\adder/norm/_0650_ ),
    .ZN(\adder/norm/_0651_ ));
 INV_X2 \adder/norm/_1556_  (.A(\adder/norm/_0651_ ),
    .ZN(\adder/norm/_0652_ ));
 NAND4_X4 \adder/norm/_1557_  (.A1(\adder/norm/_0643_ ),
    .A2(\adder/norm/_0645_ ),
    .A3(\adder/norm/_0648_ ),
    .A4(\adder/norm/_0652_ ),
    .ZN(\adder/norm/_0653_ ));
 AOI21_X1 \adder/norm/_1558_  (.A(\adder/norm/_0646_ ),
    .B1(\adder/norm/_0585_ ),
    .B2(\adder/norm/_0647_ ),
    .ZN(\adder/norm/_0654_ ));
 NAND2_X4 \adder/norm/_1559_  (.A1(\adder/norm/_0653_ ),
    .A2(\adder/norm/_0654_ ),
    .ZN(\adder/norm/_0655_ ));
 NOR2_X1 \adder/norm/_1560_  (.A1(\adder/norm/_0646_ ),
    .A2(\adder/norm/_0585_ ),
    .ZN(\adder/norm/_0656_ ));
 INV_X1 \adder/norm/_1561_  (.A(\adder/norm/_0656_ ),
    .ZN(\adder/norm/_0657_ ));
 NAND4_X4 \adder/norm/_1562_  (.A1(\adder/norm/_0643_ ),
    .A2(\adder/norm/_0645_ ),
    .A3(\adder/norm/_0657_ ),
    .A4(\adder/norm/_0652_ ),
    .ZN(\adder/norm/_0658_ ));
 NAND2_X4 \adder/norm/_1563_  (.A1(\adder/norm/_0658_ ),
    .A2(\adder/norm/_0655_ ),
    .ZN(\adder/norm/_0659_ ));
 INV_X16 \adder/norm/_1564_  (.A(\adder/norm/_0659_ ),
    .ZN(\adder/norm/_0660_ ));
 BUF_X1 input4 (.A(operand_fp16_i[12]),
    .Z(net4));
 NAND2_X1 \adder/norm/_1566_  (.A1(\adder/norm/_0660_ ),
    .A2(\adder/mant_prenorm_d[31] ),
    .ZN(\adder/norm/_0662_ ));
 NAND4_X1 \adder/norm/_1567_  (.A1(\adder/norm/_0112_ ),
    .A2(\adder/norm/_0061_ ),
    .A3(\adder/norm/_0497_ ),
    .A4(\adder/norm/_0354_ ),
    .ZN(\adder/norm/_0663_ ));
 NOR3_X1 \adder/norm/_1568_  (.A1(\adder/norm/_0663_ ),
    .A2(\adder/exp_prenorm_d[1] ),
    .A3(\adder/exp_prenorm_d[0] ),
    .ZN(\adder/norm/_0664_ ));
 NOR2_X1 \adder/norm/_1569_  (.A1(\adder/exp_prenorm_d[7] ),
    .A2(\adder/exp_prenorm_d[6] ),
    .ZN(\adder/norm/_0665_ ));
 NAND4_X2 \adder/norm/_1570_  (.A1(\adder/norm/_0664_ ),
    .A2(\adder/norm/_0585_ ),
    .A3(\adder/norm/_0647_ ),
    .A4(\adder/norm/_0665_ ),
    .ZN(\adder/norm/_0666_ ));
 INV_X1 \adder/norm/_1571_  (.A(\adder/norm/_0666_ ),
    .ZN(\adder/norm/_0667_ ));
 AOI21_X1 \adder/norm/_1572_  (.A(\adder/exp_prenorm_d[0] ),
    .B1(\adder/norm/_0667_ ),
    .B2(\adder/norm/_0616_ ),
    .ZN(\adder/norm/_0668_ ));
 NAND2_X1 \adder/norm/_1573_  (.A1(\adder/norm/_0622_ ),
    .A2(\adder/norm/_0668_ ),
    .ZN(\adder/norm/_0669_ ));
 OAI21_X4 \adder/norm/_1574_  (.A(\adder/norm/_0669_ ),
    .B1(\adder/norm/Mant_leadingOne_D[0] ),
    .B2(net257),
    .ZN(\adder/norm/_0670_ ));
 BUF_X1 input3 (.A(operand_fp16_i[11]),
    .Z(net3));
 NAND2_X1 \adder/norm/_1576_  (.A1(\adder/norm/_0662_ ),
    .A2(net84),
    .ZN(\adder/norm/_0672_ ));
 INV_X32 \adder/norm/_1577_  (.A(net83),
    .ZN(\adder/norm/_0673_ ));
 BUF_X1 input2 (.A(operand_fp16_i[10]),
    .Z(net2));
 BUF_X2 input1 (.A(operand_fp16_i[0]),
    .Z(net1));
 INV_X1 \adder/norm/_1580_  (.A(\adder/mant_prenorm_d[30] ),
    .ZN(\adder/norm/_0676_ ));
 OAI21_X1 \adder/norm/_1581_  (.A(\adder/norm/_0673_ ),
    .B1(net256),
    .B2(\adder/norm/_0676_ ),
    .ZN(\adder/norm/_0677_ ));
 NAND2_X1 \adder/norm/_1582_  (.A1(\adder/norm/_0672_ ),
    .A2(\adder/norm/_0677_ ),
    .ZN(\adder/norm/_0678_ ));
 NAND2_X1 \adder/norm/_1583_  (.A1(net257),
    .A2(\adder/norm/_1464_ ),
    .ZN(\adder/norm/_0679_ ));
 OAI21_X4 \adder/norm/_1584_  (.A(\adder/norm/_0679_ ),
    .B1(\adder/norm/Mant_leadingOne_D[1] ),
    .B2(net257),
    .ZN(\adder/norm/_0680_ ));
 INV_X16 \adder/norm/_1585_  (.A(net81),
    .ZN(\adder/norm/_0681_ ));
 TAPCELL_X1 PHY_125 ();
 TAPCELL_X1 PHY_124 ();
 NAND2_X1 \adder/norm/_1588_  (.A1(\adder/norm/_0678_ ),
    .A2(\adder/norm/_0681_ ),
    .ZN(\adder/norm/_0684_ ));
 TAPCELL_X1 PHY_123 ();
 TAPCELL_X1 PHY_122 ();
 TAPCELL_X1 PHY_121 ();
 NAND3_X1 \adder/norm/_1592_  (.A1(\adder/norm/_0660_ ),
    .A2(\adder/mant_prenorm_d[33] ),
    .A3(net84),
    .ZN(\adder/norm/_0688_ ));
 TAPCELL_X1 PHY_120 ();
 TAPCELL_X1 PHY_119 ();
 NAND3_X1 \adder/norm/_1595_  (.A1(\adder/norm/_0660_ ),
    .A2(\adder/mant_prenorm_d[32] ),
    .A3(\adder/norm/_0673_ ),
    .ZN(\adder/norm/_0691_ ));
 TAPCELL_X1 PHY_118 ();
 NAND3_X1 \adder/norm/_1597_  (.A1(\adder/norm/_0688_ ),
    .A2(\adder/norm/_0691_ ),
    .A3(net82),
    .ZN(\adder/norm/_0693_ ));
 INV_X16 \adder/norm/_1598_  (.A(net259),
    .ZN(\adder/norm/_0694_ ));
 TAPCELL_X1 PHY_117 ();
 NAND3_X1 \adder/norm/_1600_  (.A1(\adder/norm/_0684_ ),
    .A2(\adder/norm/_0693_ ),
    .A3(\adder/norm/_0694_ ),
    .ZN(\adder/norm/_0696_ ));
 TAPCELL_X1 PHY_116 ();
 NAND2_X1 \adder/norm/_1602_  (.A1(\adder/norm/_0660_ ),
    .A2(\adder/mant_prenorm_d[28] ),
    .ZN(\adder/norm/_0698_ ));
 NAND2_X1 \adder/norm/_1603_  (.A1(\adder/norm/_0698_ ),
    .A2(\adder/norm/_0673_ ),
    .ZN(\adder/norm/_0699_ ));
 TAPCELL_X1 PHY_115 ();
 INV_X1 \adder/norm/_1605_  (.A(\adder/mant_prenorm_d[29] ),
    .ZN(\adder/norm/_0701_ ));
 OAI21_X1 \adder/norm/_1606_  (.A(net84),
    .B1(\adder/norm/_0659_ ),
    .B2(\adder/norm/_0701_ ),
    .ZN(\adder/norm/_0702_ ));
 NAND2_X1 \adder/norm/_1607_  (.A1(\adder/norm/_0699_ ),
    .A2(\adder/norm/_0702_ ),
    .ZN(\adder/norm/_0703_ ));
 TAPCELL_X1 PHY_114 ();
 NAND2_X1 \adder/norm/_1609_  (.A1(\adder/norm/_0703_ ),
    .A2(net82),
    .ZN(\adder/norm/_0705_ ));
 TAPCELL_X1 PHY_113 ();
 TAPCELL_X1 PHY_112 ();
 TAPCELL_X1 PHY_111 ();
 NAND4_X1 \adder/norm/_1613_  (.A1(\adder/norm/_0655_ ),
    .A2(\adder/mant_prenorm_d[27] ),
    .A3(net84),
    .A4(net249),
    .ZN(\adder/norm/_0709_ ));
 NAND4_X1 \adder/norm/_1614_  (.A1(\adder/norm/_0655_ ),
    .A2(\adder/mant_prenorm_d[26] ),
    .A3(\adder/norm/_0673_ ),
    .A4(net249),
    .ZN(\adder/norm/_0710_ ));
 TAPCELL_X1 PHY_110 ();
 NAND3_X1 \adder/norm/_1616_  (.A1(\adder/norm/_0709_ ),
    .A2(\adder/norm/_0710_ ),
    .A3(\adder/norm/_0681_ ),
    .ZN(\adder/norm/_0712_ ));
 NAND3_X1 \adder/norm/_1617_  (.A1(\adder/norm/_0705_ ),
    .A2(net241),
    .A3(\adder/norm/_0712_ ),
    .ZN(\adder/norm/_0713_ ));
 AND2_X1 \adder/norm/_1618_  (.A1(\adder/norm/_0696_ ),
    .A2(\adder/norm/_0713_ ),
    .ZN(\adder/norm/_0714_ ));
 NAND3_X4 \adder/norm/_1619_  (.A1(net259),
    .A2(\adder/norm/_0640_ ),
    .A3(\adder/norm/_0641_ ),
    .ZN(\adder/norm/_0715_ ));
 NAND2_X4 \adder/norm/_1620_  (.A1(\adder/norm/_0694_ ),
    .A2(\adder/norm/_0642_ ),
    .ZN(\adder/norm/_0716_ ));
 NAND2_X4 \adder/norm/_1621_  (.A1(\adder/norm/_0716_ ),
    .A2(\adder/norm/_0715_ ),
    .ZN(\adder/norm/_0717_ ));
 TAPCELL_X1 PHY_109 ();
 TAPCELL_X1 PHY_108 ();
 NAND2_X1 \adder/norm/_1624_  (.A1(\adder/norm/_0714_ ),
    .A2(net250),
    .ZN(\adder/norm/_0720_ ));
 TAPCELL_X1 PHY_107 ();
 INV_X1 \adder/norm/_1626_  (.A(\adder/mant_prenorm_d[20] ),
    .ZN(\adder/norm/_0722_ ));
 OAI21_X1 \adder/norm/_1627_  (.A(\adder/norm/_0673_ ),
    .B1(\adder/norm/_0659_ ),
    .B2(\adder/norm/_0722_ ),
    .ZN(\adder/norm/_0723_ ));
 TAPCELL_X1 PHY_106 ();
 INV_X1 \adder/norm/_1629_  (.A(\adder/mant_prenorm_d[21] ),
    .ZN(\adder/norm/_0725_ ));
 OAI21_X1 \adder/norm/_1630_  (.A(net84),
    .B1(\adder/norm/_0659_ ),
    .B2(\adder/norm/_0725_ ),
    .ZN(\adder/norm/_0726_ ));
 NAND2_X1 \adder/norm/_1631_  (.A1(\adder/norm/_0723_ ),
    .A2(\adder/norm/_0726_ ),
    .ZN(\adder/norm/_0727_ ));
 NAND2_X1 \adder/norm/_1632_  (.A1(\adder/norm/_0727_ ),
    .A2(net82),
    .ZN(\adder/norm/_0728_ ));
 TAPCELL_X1 PHY_105 ();
 NAND4_X1 \adder/norm/_1634_  (.A1(\adder/norm/_0655_ ),
    .A2(net125),
    .A3(net83),
    .A4(net244),
    .ZN(\adder/norm/_0730_ ));
 NAND4_X1 \adder/norm/_1635_  (.A1(\adder/norm/_0655_ ),
    .A2(net126),
    .A3(\adder/norm/_0673_ ),
    .A4(net244),
    .ZN(\adder/norm/_0731_ ));
 NAND3_X1 \adder/norm/_1636_  (.A1(\adder/norm/_0730_ ),
    .A2(\adder/norm/_0731_ ),
    .A3(\adder/norm/_0681_ ),
    .ZN(\adder/norm/_0732_ ));
 NAND2_X1 \adder/norm/_1637_  (.A1(\adder/norm/_0728_ ),
    .A2(\adder/norm/_0732_ ),
    .ZN(\adder/norm/_0733_ ));
 TAPCELL_X1 PHY_104 ();
 NAND2_X1 \adder/norm/_1639_  (.A1(\adder/norm/_0733_ ),
    .A2(net240),
    .ZN(\adder/norm/_0735_ ));
 TAPCELL_X1 PHY_103 ();
 NAND3_X1 \adder/norm/_1641_  (.A1(\adder/norm/_0660_ ),
    .A2(\adder/mant_prenorm_d[23] ),
    .A3(net84),
    .ZN(\adder/norm/_0737_ ));
 NAND4_X1 \adder/norm/_1642_  (.A1(\adder/norm/_0655_ ),
    .A2(\adder/mant_prenorm_d[22] ),
    .A3(\adder/norm/_0673_ ),
    .A4(net268),
    .ZN(\adder/norm/_0738_ ));
 NAND3_X1 \adder/norm/_1643_  (.A1(\adder/norm/_0737_ ),
    .A2(\adder/norm/_0681_ ),
    .A3(\adder/norm/_0738_ ),
    .ZN(\adder/norm/_0739_ ));
 NAND3_X1 \adder/norm/_1644_  (.A1(\adder/norm/_0660_ ),
    .A2(\adder/mant_prenorm_d[25] ),
    .A3(net84),
    .ZN(\adder/norm/_0740_ ));
 NAND4_X1 \adder/norm/_1645_  (.A1(\adder/norm/_0655_ ),
    .A2(\adder/mant_prenorm_d[24] ),
    .A3(\adder/norm/_0673_ ),
    .A4(net268),
    .ZN(\adder/norm/_0741_ ));
 NAND3_X1 \adder/norm/_1646_  (.A1(\adder/norm/_0740_ ),
    .A2(net82),
    .A3(\adder/norm/_0741_ ),
    .ZN(\adder/norm/_0742_ ));
 NAND2_X1 \adder/norm/_1647_  (.A1(\adder/norm/_0739_ ),
    .A2(\adder/norm/_0742_ ),
    .ZN(\adder/norm/_0743_ ));
 TAPCELL_X1 PHY_102 ();
 NAND2_X1 \adder/norm/_1649_  (.A1(\adder/norm/_0743_ ),
    .A2(\adder/norm/_0694_ ),
    .ZN(\adder/norm/_0745_ ));
 NAND2_X1 \adder/norm/_1650_  (.A1(\adder/norm/_0735_ ),
    .A2(\adder/norm/_0745_ ),
    .ZN(\adder/norm/_0746_ ));
 INV_X16 \adder/norm/_1651_  (.A(\adder/norm/_0717_ ),
    .ZN(\adder/norm/_0747_ ));
 TAPCELL_X1 PHY_101 ();
 TAPCELL_X1 PHY_100 ();
 NAND2_X1 \adder/norm/_1654_  (.A1(\adder/norm/_0746_ ),
    .A2(\adder/norm/_0747_ ),
    .ZN(\adder/norm/_0750_ ));
 AND2_X2 \adder/norm/_1655_  (.A1(\adder/norm/_0643_ ),
    .A2(\adder/norm/_0645_ ),
    .ZN(\adder/norm/_0751_ ));
 INV_X1 \adder/norm/_1656_  (.A(\adder/norm/_0751_ ),
    .ZN(\adder/norm/_0752_ ));
 OR2_X1 \adder/norm/_1657_  (.A1(\adder/norm/_0643_ ),
    .A2(\adder/norm/_0645_ ),
    .ZN(\adder/norm/_0753_ ));
 NAND2_X4 \adder/norm/_1658_  (.A1(\adder/norm/_0752_ ),
    .A2(\adder/norm/_0753_ ),
    .ZN(\adder/norm/_0754_ ));
 INV_X1 \adder/norm/_1659_  (.A(\adder/norm/_0754_ ),
    .ZN(\adder/norm/_0755_ ));
 NAND2_X1 \adder/norm/_1660_  (.A1(net259),
    .A2(\adder/norm/_0642_ ),
    .ZN(\adder/norm/_0756_ ));
 NAND3_X1 \adder/norm/_1661_  (.A1(\adder/norm/_0756_ ),
    .A2(\adder/norm/_0628_ ),
    .A3(\adder/norm/_0634_ ),
    .ZN(\adder/norm/_0757_ ));
 NAND2_X2 \adder/norm/_1662_  (.A1(\adder/norm/_0757_ ),
    .A2(\adder/norm/_0643_ ),
    .ZN(\adder/norm/_0758_ ));
 INV_X2 \adder/norm/_1663_  (.A(\adder/norm/_0758_ ),
    .ZN(\adder/norm/_0759_ ));
 NAND2_X2 \adder/norm/_1664_  (.A1(\adder/norm/_0755_ ),
    .A2(\adder/norm/_0759_ ),
    .ZN(\adder/norm/_0760_ ));
 INV_X4 \adder/norm/_1665_  (.A(\adder/norm/_0760_ ),
    .ZN(\adder/norm/_0761_ ));
 TAPCELL_X1 PHY_99 ();
 TAPCELL_X1 PHY_98 ();
 NAND3_X1 \adder/norm/_1668_  (.A1(\adder/norm/_0720_ ),
    .A2(\adder/norm/_0750_ ),
    .A3(\adder/norm/_0761_ ),
    .ZN(\adder/norm/_0764_ ));
 NAND2_X1 \adder/norm/_1669_  (.A1(\adder/norm/_0660_ ),
    .A2(net127),
    .ZN(\adder/norm/_0765_ ));
 TAPCELL_X1 PHY_97 ();
 TAPCELL_X1 PHY_96 ();
 NAND2_X1 \adder/norm/_1672_  (.A1(\adder/norm/_0765_ ),
    .A2(\adder/norm/_0673_ ),
    .ZN(\adder/norm/_0768_ ));
 TAPCELL_X1 PHY_95 ();
 INV_X1 \adder/norm/_1674_  (.A(net128),
    .ZN(\adder/norm/_0770_ ));
 OAI21_X1 \adder/norm/_1675_  (.A(net83),
    .B1(net247),
    .B2(\adder/norm/_0770_ ),
    .ZN(\adder/norm/_0771_ ));
 NAND2_X1 \adder/norm/_1676_  (.A1(\adder/norm/_0768_ ),
    .A2(\adder/norm/_0771_ ),
    .ZN(\adder/norm/_0772_ ));
 TAPCELL_X1 PHY_94 ();
 NAND2_X1 \adder/norm/_1678_  (.A1(\adder/norm/_0772_ ),
    .A2(\adder/norm/_0681_ ),
    .ZN(\adder/norm/_0774_ ));
 NAND2_X4 \adder/norm/_1679_  (.A1(\adder/norm/_0660_ ),
    .A2(net129),
    .ZN(\adder/norm/_0775_ ));
 NAND2_X1 \adder/norm/_1680_  (.A1(\adder/norm/_0775_ ),
    .A2(\adder/norm/_0673_ ),
    .ZN(\adder/norm/_0776_ ));
 INV_X1 \adder/norm/_1681_  (.A(net130),
    .ZN(\adder/norm/_0777_ ));
 OAI21_X1 \adder/norm/_1682_  (.A(net83),
    .B1(net247),
    .B2(\adder/norm/_0777_ ),
    .ZN(\adder/norm/_0778_ ));
 NAND2_X1 \adder/norm/_1683_  (.A1(\adder/norm/_0776_ ),
    .A2(\adder/norm/_0778_ ),
    .ZN(\adder/norm/_0779_ ));
 TAPCELL_X1 PHY_93 ();
 TAPCELL_X1 PHY_92 ();
 NAND2_X1 \adder/norm/_1686_  (.A1(\adder/norm/_0779_ ),
    .A2(net81),
    .ZN(\adder/norm/_0782_ ));
 NAND3_X1 \adder/norm/_1687_  (.A1(\adder/norm/_0774_ ),
    .A2(\adder/norm/_0782_ ),
    .A3(net241),
    .ZN(\adder/norm/_0783_ ));
 INV_X1 \adder/norm/_1688_  (.A(net131),
    .ZN(\adder/norm/_0784_ ));
 OAI21_X1 \adder/norm/_1689_  (.A(\adder/norm/_0673_ ),
    .B1(net247),
    .B2(\adder/norm/_0784_ ),
    .ZN(\adder/norm/_0785_ ));
 INV_X1 \adder/norm/_1690_  (.A(net132),
    .ZN(\adder/norm/_0786_ ));
 OAI21_X1 \adder/norm/_1691_  (.A(net83),
    .B1(net247),
    .B2(\adder/norm/_0786_ ),
    .ZN(\adder/norm/_0787_ ));
 NAND2_X1 \adder/norm/_1692_  (.A1(\adder/norm/_0785_ ),
    .A2(\adder/norm/_0787_ ),
    .ZN(\adder/norm/_0788_ ));
 NAND2_X1 \adder/norm/_1693_  (.A1(\adder/norm/_0788_ ),
    .A2(net81),
    .ZN(\adder/norm/_0789_ ));
 NAND3_X1 \adder/norm/_1694_  (.A1(\adder/norm/_0660_ ),
    .A2(net133),
    .A3(net83),
    .ZN(\adder/norm/_0790_ ));
 TAPCELL_X1 PHY_91 ();
 NAND3_X1 \adder/norm/_1696_  (.A1(\adder/norm/_0660_ ),
    .A2(net134),
    .A3(\adder/norm/_0673_ ),
    .ZN(\adder/norm/_0792_ ));
 NAND3_X1 \adder/norm/_1697_  (.A1(\adder/norm/_0790_ ),
    .A2(\adder/norm/_0792_ ),
    .A3(\adder/norm/_0681_ ),
    .ZN(\adder/norm/_0793_ ));
 TAPCELL_X1 PHY_90 ();
 NAND3_X1 \adder/norm/_1699_  (.A1(\adder/norm/_0789_ ),
    .A2(\adder/norm/_0793_ ),
    .A3(\adder/norm/_0694_ ),
    .ZN(\adder/norm/_0795_ ));
 NAND3_X1 \adder/norm/_1700_  (.A1(\adder/norm/_0783_ ),
    .A2(\adder/norm/_0795_ ),
    .A3(\adder/norm/_0747_ ),
    .ZN(\adder/norm/_0796_ ));
 INV_X1 \adder/norm/_1701_  (.A(net135),
    .ZN(\adder/norm/_0797_ ));
 OAI21_X1 \adder/norm/_1702_  (.A(\adder/norm/_0673_ ),
    .B1(net247),
    .B2(\adder/norm/_0797_ ),
    .ZN(\adder/norm/_0798_ ));
 INV_X1 \adder/norm/_1703_  (.A(net136),
    .ZN(\adder/norm/_0799_ ));
 OAI21_X1 \adder/norm/_1704_  (.A(net83),
    .B1(net247),
    .B2(\adder/norm/_0799_ ),
    .ZN(\adder/norm/_0800_ ));
 NAND2_X1 \adder/norm/_1705_  (.A1(\adder/norm/_0798_ ),
    .A2(\adder/norm/_0800_ ),
    .ZN(\adder/norm/_0801_ ));
 NAND2_X1 \adder/norm/_1706_  (.A1(\adder/norm/_0801_ ),
    .A2(net81),
    .ZN(\adder/norm/_0802_ ));
 NAND3_X1 \adder/norm/_1707_  (.A1(\adder/norm/_0660_ ),
    .A2(net137),
    .A3(net83),
    .ZN(\adder/norm/_0803_ ));
 TAPCELL_X1 PHY_89 ();
 TAPCELL_X1 PHY_88 ();
 NAND4_X1 \adder/norm/_1710_  (.A1(\adder/norm/_0655_ ),
    .A2(net138),
    .A3(\adder/norm/_0673_ ),
    .A4(net244),
    .ZN(\adder/norm/_0806_ ));
 NAND3_X1 \adder/norm/_1711_  (.A1(\adder/norm/_0803_ ),
    .A2(\adder/norm/_0681_ ),
    .A3(\adder/norm/_0806_ ),
    .ZN(\adder/norm/_0807_ ));
 NAND3_X1 \adder/norm/_1712_  (.A1(\adder/norm/_0802_ ),
    .A2(\adder/norm/_0807_ ),
    .A3(net241),
    .ZN(\adder/norm/_0808_ ));
 INV_X1 \adder/norm/_1713_  (.A(net139),
    .ZN(\adder/norm/_0809_ ));
 OAI21_X1 \adder/norm/_1714_  (.A(\adder/norm/_0673_ ),
    .B1(net247),
    .B2(\adder/norm/_0809_ ),
    .ZN(\adder/norm/_0810_ ));
 NAND3_X1 \adder/norm/_1715_  (.A1(\adder/norm/_0655_ ),
    .A2(net140),
    .A3(net244),
    .ZN(\adder/norm/_0811_ ));
 NAND2_X1 \adder/norm/_1716_  (.A1(\adder/norm/_0811_ ),
    .A2(net83),
    .ZN(\adder/norm/_0812_ ));
 NAND2_X1 \adder/norm/_1717_  (.A1(\adder/norm/_0810_ ),
    .A2(\adder/norm/_0812_ ),
    .ZN(\adder/norm/_0813_ ));
 NAND2_X1 \adder/norm/_1718_  (.A1(\adder/norm/_0813_ ),
    .A2(net81),
    .ZN(\adder/norm/_0814_ ));
 NAND3_X1 \adder/norm/_1719_  (.A1(\adder/norm/_0660_ ),
    .A2(net141),
    .A3(net83),
    .ZN(\adder/norm/_0815_ ));
 NAND4_X1 \adder/norm/_1720_  (.A1(\adder/norm/_0655_ ),
    .A2(net142),
    .A3(\adder/norm/_0673_ ),
    .A4(net244),
    .ZN(\adder/norm/_0816_ ));
 NAND3_X1 \adder/norm/_1721_  (.A1(\adder/norm/_0815_ ),
    .A2(\adder/norm/_0681_ ),
    .A3(\adder/norm/_0816_ ),
    .ZN(\adder/norm/_0817_ ));
 NAND3_X1 \adder/norm/_1722_  (.A1(\adder/norm/_0814_ ),
    .A2(\adder/norm/_0817_ ),
    .A3(\adder/norm/_0694_ ),
    .ZN(\adder/norm/_0818_ ));
 NAND3_X1 \adder/norm/_1723_  (.A1(\adder/norm/_0808_ ),
    .A2(\adder/norm/_0818_ ),
    .A3(net250),
    .ZN(\adder/norm/_0819_ ));
 NOR2_X4 \adder/norm/_1724_  (.A1(\adder/norm/_0754_ ),
    .A2(\adder/norm/_0759_ ),
    .ZN(\adder/norm/_0820_ ));
 TAPCELL_X1 PHY_87 ();
 TAPCELL_X1 PHY_86 ();
 NAND3_X1 \adder/norm/_1727_  (.A1(\adder/norm/_0796_ ),
    .A2(\adder/norm/_0819_ ),
    .A3(\adder/norm/_0820_ ),
    .ZN(\adder/norm/_0823_ ));
 INV_X1 \adder/norm/_1728_  (.A(\adder/mant_prenorm_d[40] ),
    .ZN(\adder/norm/_0824_ ));
 OAI21_X1 \adder/norm/_1729_  (.A(\adder/norm/_0673_ ),
    .B1(\adder/norm/_0659_ ),
    .B2(\adder/norm/_0824_ ),
    .ZN(\adder/norm/_0825_ ));
 INV_X1 \adder/norm/_1730_  (.A(\adder/mant_prenorm_d[41] ),
    .ZN(\adder/norm/_0826_ ));
 OAI21_X1 \adder/norm/_1731_  (.A(net84),
    .B1(\adder/norm/_0659_ ),
    .B2(\adder/norm/_0826_ ),
    .ZN(\adder/norm/_0827_ ));
 NAND2_X1 \adder/norm/_1732_  (.A1(\adder/norm/_0825_ ),
    .A2(\adder/norm/_0827_ ),
    .ZN(\adder/norm/_0828_ ));
 NAND2_X1 \adder/norm/_1733_  (.A1(\adder/norm/_0828_ ),
    .A2(net81),
    .ZN(\adder/norm/_0829_ ));
 TAPCELL_X1 PHY_85 ();
 TAPCELL_X1 PHY_84 ();
 TAPCELL_X1 PHY_83 ();
 TAPCELL_X1 PHY_82 ();
 NAND4_X1 \adder/norm/_1738_  (.A1(\adder/norm/_0655_ ),
    .A2(\adder/mant_prenorm_d[39] ),
    .A3(net84),
    .A4(net249),
    .ZN(\adder/norm/_0834_ ));
 NAND4_X1 \adder/norm/_1739_  (.A1(\adder/norm/_0655_ ),
    .A2(\adder/mant_prenorm_d[38] ),
    .A3(\adder/norm/_0673_ ),
    .A4(net249),
    .ZN(\adder/norm/_0835_ ));
 NAND3_X1 \adder/norm/_1740_  (.A1(\adder/norm/_0834_ ),
    .A2(\adder/norm/_0835_ ),
    .A3(\adder/norm/_0681_ ),
    .ZN(\adder/norm/_0836_ ));
 TAPCELL_X1 PHY_81 ();
 NAND3_X1 \adder/norm/_1742_  (.A1(\adder/norm/_0829_ ),
    .A2(\adder/norm/_0836_ ),
    .A3(\adder/norm/_0694_ ),
    .ZN(\adder/norm/_0838_ ));
 NAND3_X1 \adder/norm/_1743_  (.A1(\adder/norm/_0660_ ),
    .A2(\adder/mant_prenorm_d[35] ),
    .A3(net84),
    .ZN(\adder/norm/_0839_ ));
 NAND4_X1 \adder/norm/_1744_  (.A1(\adder/norm/_0655_ ),
    .A2(\adder/mant_prenorm_d[34] ),
    .A3(\adder/norm/_0673_ ),
    .A4(net268),
    .ZN(\adder/norm/_0840_ ));
 NAND3_X1 \adder/norm/_1745_  (.A1(\adder/norm/_0839_ ),
    .A2(\adder/norm/_0681_ ),
    .A3(\adder/norm/_0840_ ),
    .ZN(\adder/norm/_0841_ ));
 TAPCELL_X1 PHY_80 ();
 TAPCELL_X1 PHY_79 ();
 TAPCELL_X1 PHY_78 ();
 NAND3_X1 \adder/norm/_1749_  (.A1(\adder/norm/_0660_ ),
    .A2(\adder/mant_prenorm_d[37] ),
    .A3(net84),
    .ZN(\adder/norm/_0845_ ));
 TAPCELL_X1 PHY_77 ();
 NAND4_X1 \adder/norm/_1751_  (.A1(\adder/norm/_0655_ ),
    .A2(\adder/mant_prenorm_d[36] ),
    .A3(\adder/norm/_0673_ ),
    .A4(net249),
    .ZN(\adder/norm/_0847_ ));
 NAND3_X1 \adder/norm/_1752_  (.A1(\adder/norm/_0845_ ),
    .A2(net82),
    .A3(\adder/norm/_0847_ ),
    .ZN(\adder/norm/_0848_ ));
 TAPCELL_X1 PHY_76 ();
 NAND3_X1 \adder/norm/_1754_  (.A1(\adder/norm/_0841_ ),
    .A2(\adder/norm/_0848_ ),
    .A3(net241),
    .ZN(\adder/norm/_0850_ ));
 NAND3_X1 \adder/norm/_1755_  (.A1(\adder/norm/_0838_ ),
    .A2(\adder/norm/_0850_ ),
    .A3(\adder/norm/_0747_ ),
    .ZN(\adder/norm/_0851_ ));
 NAND3_X1 \adder/norm/_1756_  (.A1(\adder/norm/_0660_ ),
    .A2(\adder/mant_prenorm_d[45] ),
    .A3(\adder/norm/_0670_ ),
    .ZN(\adder/norm/_0852_ ));
 NAND3_X1 \adder/norm/_1757_  (.A1(\adder/norm/_0660_ ),
    .A2(\adder/mant_prenorm_d[44] ),
    .A3(\adder/norm/_0673_ ),
    .ZN(\adder/norm/_0853_ ));
 NAND3_X1 \adder/norm/_1758_  (.A1(\adder/norm/_0852_ ),
    .A2(\adder/norm/_0853_ ),
    .A3(net82),
    .ZN(\adder/norm/_0854_ ));
 NAND3_X1 \adder/norm/_1759_  (.A1(\adder/norm/_0660_ ),
    .A2(\adder/mant_prenorm_d[43] ),
    .A3(net84),
    .ZN(\adder/norm/_0855_ ));
 TAPCELL_X1 PHY_75 ();
 NAND4_X1 \adder/norm/_1761_  (.A1(\adder/norm/_0655_ ),
    .A2(\adder/mant_prenorm_d[42] ),
    .A3(\adder/norm/_0673_ ),
    .A4(net249),
    .ZN(\adder/norm/_0857_ ));
 NAND3_X1 \adder/norm/_1762_  (.A1(\adder/norm/_0855_ ),
    .A2(\adder/norm/_0681_ ),
    .A3(\adder/norm/_0857_ ),
    .ZN(\adder/norm/_0858_ ));
 TAPCELL_X1 PHY_74 ();
 NAND3_X1 \adder/norm/_1764_  (.A1(\adder/norm/_0854_ ),
    .A2(\adder/norm/_0858_ ),
    .A3(net241),
    .ZN(\adder/norm/_0860_ ));
 NAND3_X1 \adder/norm/_1765_  (.A1(\adder/norm/_0660_ ),
    .A2(\adder/mant_prenorm_d[47] ),
    .A3(net84),
    .ZN(\adder/norm/_0861_ ));
 TAPCELL_X1 PHY_73 ();
 NAND4_X1 \adder/norm/_1767_  (.A1(\adder/norm/_0655_ ),
    .A2(\adder/mant_prenorm_d[46] ),
    .A3(\adder/norm/_0673_ ),
    .A4(net249),
    .ZN(\adder/norm/_0863_ ));
 NAND2_X1 \adder/norm/_1768_  (.A1(\adder/norm/_0861_ ),
    .A2(\adder/norm/_0863_ ),
    .ZN(\adder/norm/_0864_ ));
 TAPCELL_X1 PHY_72 ();
 TAPCELL_X1 PHY_71 ();
 NAND3_X1 \adder/norm/_1771_  (.A1(\adder/norm/_0864_ ),
    .A2(\adder/norm/_0694_ ),
    .A3(\adder/norm/_0681_ ),
    .ZN(\adder/norm/_0867_ ));
 NAND3_X1 \adder/norm/_1772_  (.A1(\adder/norm/_0860_ ),
    .A2(\adder/norm/_0717_ ),
    .A3(\adder/norm/_0867_ ),
    .ZN(\adder/norm/_0868_ ));
 NAND2_X4 \adder/norm/_1773_  (.A1(\adder/norm/_0754_ ),
    .A2(\adder/norm/_0758_ ),
    .ZN(\adder/norm/_0869_ ));
 INV_X4 \adder/norm/_1774_  (.A(\adder/norm/_0869_ ),
    .ZN(\adder/norm/_0870_ ));
 TAPCELL_X1 PHY_70 ();
 NAND3_X1 \adder/norm/_1776_  (.A1(\adder/norm/_0851_ ),
    .A2(\adder/norm/_0868_ ),
    .A3(\adder/norm/_0870_ ),
    .ZN(\adder/norm/_0872_ ));
 OR2_X1 \adder/norm/_1777_  (.A1(\adder/norm/_0751_ ),
    .A2(\adder/norm/_0649_ ),
    .ZN(\adder/norm/_0873_ ));
 NAND2_X2 \adder/norm/_1778_  (.A1(\adder/norm/_0751_ ),
    .A2(\adder/norm/_0649_ ),
    .ZN(\adder/norm/_0874_ ));
 NAND2_X2 \adder/norm/_1779_  (.A1(\adder/norm/_0873_ ),
    .A2(\adder/norm/_0874_ ),
    .ZN(\adder/norm/_0875_ ));
 NAND4_X1 \adder/norm/_1780_  (.A1(\adder/norm/_0764_ ),
    .A2(\adder/norm/_0823_ ),
    .A3(\adder/norm/_0872_ ),
    .A4(\adder/norm/_0875_ ),
    .ZN(\adder/norm/_0876_ ));
 XNOR2_X2 \adder/norm/_1781_  (.A(\adder/norm/_0650_ ),
    .B(\adder/norm/_0874_ ),
    .ZN(\adder/norm/_0877_ ));
 INV_X1 \adder/norm/_1782_  (.A(net143),
    .ZN(\adder/norm/_0878_ ));
 OAI21_X1 \adder/norm/_1783_  (.A(\adder/norm/_0673_ ),
    .B1(net247),
    .B2(\adder/norm/_0878_ ),
    .ZN(\adder/norm/_0879_ ));
 TAPCELL_X1 PHY_69 ();
 NAND3_X1 \adder/norm/_1785_  (.A1(\adder/norm/_0655_ ),
    .A2(net144),
    .A3(net244),
    .ZN(\adder/norm/_0881_ ));
 NAND2_X1 \adder/norm/_1786_  (.A1(\adder/norm/_0881_ ),
    .A2(net83),
    .ZN(\adder/norm/_0882_ ));
 NAND3_X1 \adder/norm/_1787_  (.A1(\adder/norm/_0879_ ),
    .A2(net81),
    .A3(\adder/norm/_0882_ ),
    .ZN(\adder/norm/_0883_ ));
 TAPCELL_X1 PHY_68 ();
 NOR2_X1 \adder/norm/_1789_  (.A1(\adder/norm/_0883_ ),
    .A2(net240),
    .ZN(\adder/norm/_0885_ ));
 INV_X1 \adder/norm/_1790_  (.A(\adder/norm/_0885_ ),
    .ZN(\adder/norm/_0886_ ));
 NOR2_X1 \adder/norm/_1791_  (.A1(\adder/norm/_0886_ ),
    .A2(\adder/norm/_0747_ ),
    .ZN(\adder/norm/_0887_ ));
 NAND2_X4 \adder/norm/_1792_  (.A1(\adder/norm/_0754_ ),
    .A2(\adder/norm/_0759_ ),
    .ZN(\adder/norm/_0888_ ));
 INV_X4 \adder/norm/_1793_  (.A(\adder/norm/_0888_ ),
    .ZN(\adder/norm/_0889_ ));
 TAPCELL_X1 PHY_67 ();
 NAND2_X1 \adder/norm/_1795_  (.A1(\adder/norm/_0887_ ),
    .A2(\adder/norm/_0889_ ),
    .ZN(\adder/norm/_0891_ ));
 INV_X4 \adder/norm/_1796_  (.A(\adder/norm/_0875_ ),
    .ZN(\adder/norm/_0892_ ));
 TAPCELL_X1 PHY_66 ();
 TAPCELL_X1 PHY_65 ();
 AOI21_X1 \adder/norm/_1799_  (.A(\adder/norm/_0877_ ),
    .B1(\adder/norm/_0891_ ),
    .B2(\adder/norm/_0892_ ),
    .ZN(\adder/norm/_0895_ ));
 NAND2_X1 \adder/norm/_1800_  (.A1(\adder/norm/_0876_ ),
    .A2(\adder/norm/_0895_ ),
    .ZN(\adder/norm/_0896_ ));
 NAND2_X1 \adder/norm/_1801_  (.A1(\adder/norm/_0660_ ),
    .A2(\adder/mant_prenorm_d[23] ),
    .ZN(\adder/norm/_0897_ ));
 NAND2_X1 \adder/norm/_1802_  (.A1(\adder/norm/_0897_ ),
    .A2(\adder/norm/_0673_ ),
    .ZN(\adder/norm/_0898_ ));
 NAND2_X1 \adder/norm/_1803_  (.A1(\adder/norm/_0660_ ),
    .A2(\adder/mant_prenorm_d[24] ),
    .ZN(\adder/norm/_0899_ ));
 NAND2_X1 \adder/norm/_1804_  (.A1(\adder/norm/_0899_ ),
    .A2(net83),
    .ZN(\adder/norm/_0900_ ));
 NAND2_X1 \adder/norm/_1805_  (.A1(\adder/norm/_0898_ ),
    .A2(\adder/norm/_0900_ ),
    .ZN(\adder/norm/_0901_ ));
 NAND2_X1 \adder/norm/_1806_  (.A1(\adder/norm/_0901_ ),
    .A2(net81),
    .ZN(\adder/norm/_0902_ ));
 NAND3_X1 \adder/norm/_1807_  (.A1(\adder/norm/_0660_ ),
    .A2(\adder/mant_prenorm_d[22] ),
    .A3(net83),
    .ZN(\adder/norm/_0903_ ));
 NAND4_X1 \adder/norm/_1808_  (.A1(\adder/norm/_0655_ ),
    .A2(\adder/mant_prenorm_d[21] ),
    .A3(\adder/norm/_0673_ ),
    .A4(net249),
    .ZN(\adder/norm/_0904_ ));
 NAND3_X1 \adder/norm/_1809_  (.A1(\adder/norm/_0903_ ),
    .A2(\adder/norm/_0681_ ),
    .A3(\adder/norm/_0904_ ),
    .ZN(\adder/norm/_0905_ ));
 NAND2_X1 \adder/norm/_1810_  (.A1(\adder/norm/_0902_ ),
    .A2(\adder/norm/_0905_ ),
    .ZN(\adder/norm/_0906_ ));
 TAPCELL_X1 PHY_64 ();
 NAND2_X1 \adder/norm/_1812_  (.A1(\adder/norm/_0906_ ),
    .A2(\adder/norm/_0694_ ),
    .ZN(\adder/norm/_0908_ ));
 NAND3_X1 \adder/norm/_1813_  (.A1(\adder/norm/_0660_ ),
    .A2(\adder/mant_prenorm_d[20] ),
    .A3(net83),
    .ZN(\adder/norm/_0909_ ));
 NAND3_X1 \adder/norm/_1814_  (.A1(\adder/norm/_0660_ ),
    .A2(net145),
    .A3(\adder/norm/_0673_ ),
    .ZN(\adder/norm/_0910_ ));
 NAND3_X1 \adder/norm/_1815_  (.A1(\adder/norm/_0909_ ),
    .A2(\adder/norm/_0910_ ),
    .A3(net81),
    .ZN(\adder/norm/_0911_ ));
 NAND4_X1 \adder/norm/_1816_  (.A1(\adder/norm/_0655_ ),
    .A2(net146),
    .A3(net83),
    .A4(net244),
    .ZN(\adder/norm/_0912_ ));
 NAND4_X1 \adder/norm/_1817_  (.A1(\adder/norm/_0655_ ),
    .A2(net147),
    .A3(\adder/norm/_0673_ ),
    .A4(net244),
    .ZN(\adder/norm/_0913_ ));
 NAND3_X1 \adder/norm/_1818_  (.A1(\adder/norm/_0912_ ),
    .A2(\adder/norm/_0913_ ),
    .A3(\adder/norm/_0681_ ),
    .ZN(\adder/norm/_0914_ ));
 NAND2_X1 \adder/norm/_1819_  (.A1(\adder/norm/_0911_ ),
    .A2(\adder/norm/_0914_ ),
    .ZN(\adder/norm/_0915_ ));
 NAND2_X1 \adder/norm/_1820_  (.A1(\adder/norm/_0915_ ),
    .A2(net240),
    .ZN(\adder/norm/_0916_ ));
 NAND2_X1 \adder/norm/_1821_  (.A1(\adder/norm/_0908_ ),
    .A2(\adder/norm/_0916_ ),
    .ZN(\adder/norm/_0917_ ));
 NAND2_X1 \adder/norm/_1822_  (.A1(\adder/norm/_0917_ ),
    .A2(\adder/norm/_0747_ ),
    .ZN(\adder/norm/_0918_ ));
 INV_X1 \adder/norm/_1823_  (.A(\adder/mant_prenorm_d[26] ),
    .ZN(\adder/norm/_0919_ ));
 OAI21_X1 \adder/norm/_1824_  (.A(net84),
    .B1(net256),
    .B2(\adder/norm/_0919_ ),
    .ZN(\adder/norm/_0920_ ));
 INV_X1 \adder/norm/_1825_  (.A(\adder/mant_prenorm_d[25] ),
    .ZN(\adder/norm/_0921_ ));
 OAI21_X1 \adder/norm/_1826_  (.A(\adder/norm/_0673_ ),
    .B1(net256),
    .B2(\adder/norm/_0921_ ),
    .ZN(\adder/norm/_0922_ ));
 NAND2_X1 \adder/norm/_1827_  (.A1(\adder/norm/_0920_ ),
    .A2(\adder/norm/_0922_ ),
    .ZN(\adder/norm/_0923_ ));
 NAND2_X1 \adder/norm/_1828_  (.A1(\adder/norm/_0923_ ),
    .A2(\adder/norm/_0681_ ),
    .ZN(\adder/norm/_0924_ ));
 NAND3_X1 \adder/norm/_1829_  (.A1(\adder/norm/_0660_ ),
    .A2(\adder/mant_prenorm_d[28] ),
    .A3(net83),
    .ZN(\adder/norm/_0925_ ));
 NAND3_X1 \adder/norm/_1830_  (.A1(\adder/norm/_0660_ ),
    .A2(\adder/mant_prenorm_d[27] ),
    .A3(\adder/norm/_0673_ ),
    .ZN(\adder/norm/_0926_ ));
 NAND3_X1 \adder/norm/_1831_  (.A1(\adder/norm/_0925_ ),
    .A2(\adder/norm/_0926_ ),
    .A3(net81),
    .ZN(\adder/norm/_0927_ ));
 NAND3_X1 \adder/norm/_1832_  (.A1(\adder/norm/_0924_ ),
    .A2(\adder/norm/_0927_ ),
    .A3(net241),
    .ZN(\adder/norm/_0928_ ));
 NAND3_X1 \adder/norm/_1833_  (.A1(\adder/norm/_0660_ ),
    .A2(\adder/mant_prenorm_d[32] ),
    .A3(net83),
    .ZN(\adder/norm/_0929_ ));
 NAND3_X1 \adder/norm/_1834_  (.A1(\adder/norm/_0660_ ),
    .A2(\adder/mant_prenorm_d[31] ),
    .A3(\adder/norm/_0673_ ),
    .ZN(\adder/norm/_0930_ ));
 NAND3_X1 \adder/norm/_1835_  (.A1(\adder/norm/_0929_ ),
    .A2(\adder/norm/_0930_ ),
    .A3(net81),
    .ZN(\adder/norm/_0931_ ));
 NAND3_X1 \adder/norm/_1836_  (.A1(\adder/norm/_0660_ ),
    .A2(\adder/mant_prenorm_d[30] ),
    .A3(net83),
    .ZN(\adder/norm/_0932_ ));
 NAND4_X1 \adder/norm/_1837_  (.A1(\adder/norm/_0655_ ),
    .A2(\adder/mant_prenorm_d[29] ),
    .A3(\adder/norm/_0673_ ),
    .A4(net268),
    .ZN(\adder/norm/_0933_ ));
 NAND3_X1 \adder/norm/_1838_  (.A1(\adder/norm/_0932_ ),
    .A2(\adder/norm/_0681_ ),
    .A3(\adder/norm/_0933_ ),
    .ZN(\adder/norm/_0934_ ));
 NAND3_X1 \adder/norm/_1839_  (.A1(\adder/norm/_0931_ ),
    .A2(\adder/norm/_0934_ ),
    .A3(\adder/norm/_0694_ ),
    .ZN(\adder/norm/_0935_ ));
 NAND3_X1 \adder/norm/_1840_  (.A1(\adder/norm/_0928_ ),
    .A2(\adder/norm/_0935_ ),
    .A3(net250),
    .ZN(\adder/norm/_0936_ ));
 NAND3_X1 \adder/norm/_1841_  (.A1(\adder/norm/_0918_ ),
    .A2(\adder/norm/_0936_ ),
    .A3(\adder/norm/_0761_ ),
    .ZN(\adder/norm/_0937_ ));
 NAND2_X1 \adder/norm/_1842_  (.A1(\adder/norm/_0775_ ),
    .A2(net83),
    .ZN(\adder/norm/_0938_ ));
 OAI21_X1 \adder/norm/_1843_  (.A(\adder/norm/_0673_ ),
    .B1(net247),
    .B2(\adder/norm/_0770_ ),
    .ZN(\adder/norm/_0939_ ));
 NAND2_X1 \adder/norm/_1844_  (.A1(\adder/norm/_0938_ ),
    .A2(\adder/norm/_0939_ ),
    .ZN(\adder/norm/_0940_ ));
 NAND2_X1 \adder/norm/_1845_  (.A1(\adder/norm/_0940_ ),
    .A2(net81),
    .ZN(\adder/norm/_0941_ ));
 NAND3_X4 \adder/norm/_1846_  (.A1(\adder/norm/_0660_ ),
    .A2(net148),
    .A3(net258),
    .ZN(\adder/norm/_0942_ ));
 NAND4_X1 \adder/norm/_1847_  (.A1(\adder/norm/_0655_ ),
    .A2(net149),
    .A3(\adder/norm/_0673_ ),
    .A4(net244),
    .ZN(\adder/norm/_0943_ ));
 NAND3_X1 \adder/norm/_1848_  (.A1(\adder/norm/_0942_ ),
    .A2(\adder/norm/_0681_ ),
    .A3(\adder/norm/_0943_ ),
    .ZN(\adder/norm/_0944_ ));
 NAND3_X1 \adder/norm/_1849_  (.A1(\adder/norm/_0941_ ),
    .A2(\adder/norm/_0944_ ),
    .A3(net241),
    .ZN(\adder/norm/_0945_ ));
 NAND3_X2 \adder/norm/_1850_  (.A1(\adder/norm/_0660_ ),
    .A2(net150),
    .A3(net258),
    .ZN(\adder/norm/_0946_ ));
 NAND4_X1 \adder/norm/_1851_  (.A1(\adder/norm/_0655_ ),
    .A2(net151),
    .A3(\adder/norm/_0673_ ),
    .A4(net244),
    .ZN(\adder/norm/_0947_ ));
 NAND3_X1 \adder/norm/_1852_  (.A1(\adder/norm/_0946_ ),
    .A2(\adder/norm/_0681_ ),
    .A3(\adder/norm/_0947_ ),
    .ZN(\adder/norm/_0948_ ));
 NAND3_X2 \adder/norm/_1853_  (.A1(\adder/norm/_0660_ ),
    .A2(net152),
    .A3(net258),
    .ZN(\adder/norm/_0949_ ));
 NAND4_X1 \adder/norm/_1854_  (.A1(\adder/norm/_0655_ ),
    .A2(net153),
    .A3(\adder/norm/_0673_ ),
    .A4(net244),
    .ZN(\adder/norm/_0950_ ));
 NAND3_X1 \adder/norm/_1855_  (.A1(\adder/norm/_0949_ ),
    .A2(net81),
    .A3(\adder/norm/_0950_ ),
    .ZN(\adder/norm/_0951_ ));
 NAND3_X1 \adder/norm/_1856_  (.A1(\adder/norm/_0948_ ),
    .A2(\adder/norm/_0951_ ),
    .A3(\adder/norm/_0694_ ),
    .ZN(\adder/norm/_0952_ ));
 NAND3_X1 \adder/norm/_1857_  (.A1(\adder/norm/_0945_ ),
    .A2(\adder/norm/_0952_ ),
    .A3(\adder/norm/_0747_ ),
    .ZN(\adder/norm/_0953_ ));
 NAND3_X1 \adder/norm/_1858_  (.A1(\adder/norm/_0660_ ),
    .A2(net154),
    .A3(net83),
    .ZN(\adder/norm/_0954_ ));
 NAND4_X1 \adder/norm/_1859_  (.A1(\adder/norm/_0655_ ),
    .A2(net155),
    .A3(\adder/norm/_0673_ ),
    .A4(net244),
    .ZN(\adder/norm/_0955_ ));
 NAND3_X1 \adder/norm/_1860_  (.A1(\adder/norm/_0954_ ),
    .A2(net81),
    .A3(\adder/norm/_0955_ ),
    .ZN(\adder/norm/_0956_ ));
 NAND4_X1 \adder/norm/_1861_  (.A1(\adder/norm/_0655_ ),
    .A2(net156),
    .A3(net258),
    .A4(net244),
    .ZN(\adder/norm/_0957_ ));
 NAND4_X1 \adder/norm/_1862_  (.A1(\adder/norm/_0655_ ),
    .A2(net157),
    .A3(\adder/norm/_0673_ ),
    .A4(net244),
    .ZN(\adder/norm/_0958_ ));
 NAND3_X1 \adder/norm/_1863_  (.A1(\adder/norm/_0957_ ),
    .A2(\adder/norm/_0958_ ),
    .A3(\adder/norm/_0681_ ),
    .ZN(\adder/norm/_0959_ ));
 NAND2_X1 \adder/norm/_1864_  (.A1(\adder/norm/_0956_ ),
    .A2(\adder/norm/_0959_ ),
    .ZN(\adder/norm/_0960_ ));
 NAND2_X1 \adder/norm/_1865_  (.A1(\adder/norm/_0960_ ),
    .A2(net240),
    .ZN(\adder/norm/_0961_ ));
 NAND4_X1 \adder/norm/_1866_  (.A1(\adder/norm/_0655_ ),
    .A2(net158),
    .A3(net83),
    .A4(net244),
    .ZN(\adder/norm/_0962_ ));
 NAND4_X1 \adder/norm/_1867_  (.A1(\adder/norm/_0655_ ),
    .A2(net159),
    .A3(\adder/norm/_0673_ ),
    .A4(net244),
    .ZN(\adder/norm/_0963_ ));
 NAND3_X1 \adder/norm/_1868_  (.A1(\adder/norm/_0962_ ),
    .A2(\adder/norm/_0963_ ),
    .A3(\adder/norm/_0681_ ),
    .ZN(\adder/norm/_0964_ ));
 NAND4_X1 \adder/norm/_1869_  (.A1(\adder/norm/_0655_ ),
    .A2(net160),
    .A3(net83),
    .A4(net244),
    .ZN(\adder/norm/_0965_ ));
 NAND4_X1 \adder/norm/_1870_  (.A1(\adder/norm/_0655_ ),
    .A2(net161),
    .A3(\adder/norm/_0673_ ),
    .A4(net244),
    .ZN(\adder/norm/_0966_ ));
 NAND3_X1 \adder/norm/_1871_  (.A1(\adder/norm/_0965_ ),
    .A2(\adder/norm/_0966_ ),
    .A3(net81),
    .ZN(\adder/norm/_0967_ ));
 NAND2_X1 \adder/norm/_1872_  (.A1(\adder/norm/_0964_ ),
    .A2(\adder/norm/_0967_ ),
    .ZN(\adder/norm/_0968_ ));
 NAND2_X1 \adder/norm/_1873_  (.A1(\adder/norm/_0968_ ),
    .A2(\adder/norm/_0694_ ),
    .ZN(\adder/norm/_0969_ ));
 NAND2_X1 \adder/norm/_1874_  (.A1(\adder/norm/_0961_ ),
    .A2(\adder/norm/_0969_ ),
    .ZN(\adder/norm/_0970_ ));
 NAND2_X1 \adder/norm/_1875_  (.A1(\adder/norm/_0970_ ),
    .A2(net250),
    .ZN(\adder/norm/_0971_ ));
 NAND3_X1 \adder/norm/_1876_  (.A1(\adder/norm/_0953_ ),
    .A2(\adder/norm/_0971_ ),
    .A3(\adder/norm/_0820_ ),
    .ZN(\adder/norm/_0972_ ));
 NAND3_X1 \adder/norm/_1877_  (.A1(\adder/norm/_0660_ ),
    .A2(\adder/mant_prenorm_d[34] ),
    .A3(net83),
    .ZN(\adder/norm/_0973_ ));
 NAND4_X1 \adder/norm/_1878_  (.A1(\adder/norm/_0655_ ),
    .A2(\adder/mant_prenorm_d[33] ),
    .A3(\adder/norm/_0673_ ),
    .A4(net268),
    .ZN(\adder/norm/_0974_ ));
 NAND3_X1 \adder/norm/_1879_  (.A1(\adder/norm/_0973_ ),
    .A2(\adder/norm/_0681_ ),
    .A3(\adder/norm/_0974_ ),
    .ZN(\adder/norm/_0975_ ));
 NAND3_X1 \adder/norm/_1880_  (.A1(\adder/norm/_0660_ ),
    .A2(\adder/mant_prenorm_d[36] ),
    .A3(net84),
    .ZN(\adder/norm/_0976_ ));
 NAND4_X1 \adder/norm/_1881_  (.A1(\adder/norm/_0655_ ),
    .A2(\adder/mant_prenorm_d[35] ),
    .A3(\adder/norm/_0673_ ),
    .A4(net268),
    .ZN(\adder/norm/_0977_ ));
 NAND3_X1 \adder/norm/_1882_  (.A1(\adder/norm/_0976_ ),
    .A2(net82),
    .A3(\adder/norm/_0977_ ),
    .ZN(\adder/norm/_0978_ ));
 NAND3_X1 \adder/norm/_1883_  (.A1(\adder/norm/_0975_ ),
    .A2(\adder/norm/_0978_ ),
    .A3(net241),
    .ZN(\adder/norm/_0979_ ));
 NAND3_X1 \adder/norm/_1884_  (.A1(\adder/norm/_0660_ ),
    .A2(\adder/mant_prenorm_d[40] ),
    .A3(\adder/norm/_0670_ ),
    .ZN(\adder/norm/_0980_ ));
 NAND4_X1 \adder/norm/_1885_  (.A1(\adder/norm/_0655_ ),
    .A2(\adder/mant_prenorm_d[39] ),
    .A3(\adder/norm/_0673_ ),
    .A4(\adder/norm/_0658_ ),
    .ZN(\adder/norm/_0981_ ));
 NAND3_X1 \adder/norm/_1886_  (.A1(\adder/norm/_0980_ ),
    .A2(\adder/norm/_0680_ ),
    .A3(\adder/norm/_0981_ ),
    .ZN(\adder/norm/_0982_ ));
 NAND4_X1 \adder/norm/_1887_  (.A1(\adder/norm/_0655_ ),
    .A2(\adder/mant_prenorm_d[38] ),
    .A3(\adder/norm/_0670_ ),
    .A4(net249),
    .ZN(\adder/norm/_0983_ ));
 NAND4_X1 \adder/norm/_1888_  (.A1(\adder/norm/_0655_ ),
    .A2(\adder/mant_prenorm_d[37] ),
    .A3(\adder/norm/_0673_ ),
    .A4(\adder/norm/_0658_ ),
    .ZN(\adder/norm/_0984_ ));
 NAND3_X1 \adder/norm/_1889_  (.A1(\adder/norm/_0983_ ),
    .A2(\adder/norm/_0984_ ),
    .A3(\adder/norm/_0681_ ),
    .ZN(\adder/norm/_0985_ ));
 NAND3_X1 \adder/norm/_1890_  (.A1(\adder/norm/_0982_ ),
    .A2(\adder/norm/_0985_ ),
    .A3(\adder/norm/_0694_ ),
    .ZN(\adder/norm/_0986_ ));
 TAPCELL_X1 PHY_63 ();
 TAPCELL_X1 PHY_62 ();
 NAND3_X1 \adder/norm/_1893_  (.A1(\adder/norm/_0979_ ),
    .A2(\adder/norm/_0986_ ),
    .A3(\adder/norm/_0747_ ),
    .ZN(\adder/norm/_0989_ ));
 NAND3_X1 \adder/norm/_1894_  (.A1(\adder/norm/_0660_ ),
    .A2(\adder/mant_prenorm_d[44] ),
    .A3(net258),
    .ZN(\adder/norm/_0990_ ));
 NAND4_X1 \adder/norm/_1895_  (.A1(\adder/norm/_0655_ ),
    .A2(\adder/mant_prenorm_d[43] ),
    .A3(\adder/norm/_0673_ ),
    .A4(\adder/norm/_0658_ ),
    .ZN(\adder/norm/_0991_ ));
 NAND3_X1 \adder/norm/_1896_  (.A1(\adder/norm/_0990_ ),
    .A2(\adder/norm/_0680_ ),
    .A3(\adder/norm/_0991_ ),
    .ZN(\adder/norm/_0992_ ));
 NAND4_X1 \adder/norm/_1897_  (.A1(\adder/norm/_0655_ ),
    .A2(\adder/mant_prenorm_d[42] ),
    .A3(\adder/norm/_0670_ ),
    .A4(net249),
    .ZN(\adder/norm/_0993_ ));
 NAND4_X1 \adder/norm/_1898_  (.A1(\adder/norm/_0655_ ),
    .A2(\adder/mant_prenorm_d[41] ),
    .A3(\adder/norm/_0673_ ),
    .A4(net249),
    .ZN(\adder/norm/_0994_ ));
 NAND3_X1 \adder/norm/_1899_  (.A1(\adder/norm/_0993_ ),
    .A2(\adder/norm/_0994_ ),
    .A3(\adder/norm/_0681_ ),
    .ZN(\adder/norm/_0995_ ));
 NAND3_X1 \adder/norm/_1900_  (.A1(\adder/norm/_0992_ ),
    .A2(\adder/norm/_0995_ ),
    .A3(net241),
    .ZN(\adder/norm/_0996_ ));
 NAND4_X1 \adder/norm/_1901_  (.A1(\adder/norm/_0655_ ),
    .A2(\adder/mant_prenorm_d[46] ),
    .A3(net258),
    .A4(net244),
    .ZN(\adder/norm/_0997_ ));
 NAND4_X1 \adder/norm/_1902_  (.A1(\adder/norm/_0655_ ),
    .A2(\adder/mant_prenorm_d[45] ),
    .A3(\adder/norm/_0673_ ),
    .A4(net244),
    .ZN(\adder/norm/_0998_ ));
 NAND3_X1 \adder/norm/_1903_  (.A1(\adder/norm/_0997_ ),
    .A2(\adder/norm/_0998_ ),
    .A3(\adder/norm/_0681_ ),
    .ZN(\adder/norm/_0999_ ));
 NAND3_X1 \adder/norm/_1904_  (.A1(\adder/norm/_0660_ ),
    .A2(\adder/mant_prenorm_d[47] ),
    .A3(\adder/norm/_0673_ ),
    .ZN(\adder/norm/_1000_ ));
 NAND2_X1 \adder/norm/_1905_  (.A1(\adder/norm/_1000_ ),
    .A2(\adder/norm/_0680_ ),
    .ZN(\adder/norm/_1001_ ));
 NAND3_X1 \adder/norm/_1906_  (.A1(\adder/norm/_0999_ ),
    .A2(\adder/norm/_1001_ ),
    .A3(\adder/norm/_0694_ ),
    .ZN(\adder/norm/_1002_ ));
 TAPCELL_X1 PHY_61 ();
 TAPCELL_X1 PHY_60 ();
 NAND3_X1 \adder/norm/_1909_  (.A1(\adder/norm/_0996_ ),
    .A2(\adder/norm/_1002_ ),
    .A3(\adder/norm/_0717_ ),
    .ZN(\adder/norm/_1005_ ));
 NAND3_X1 \adder/norm/_1910_  (.A1(\adder/norm/_0989_ ),
    .A2(\adder/norm/_1005_ ),
    .A3(\adder/norm/_0870_ ),
    .ZN(\adder/norm/_1006_ ));
 NAND4_X1 \adder/norm/_1911_  (.A1(\adder/norm/_0937_ ),
    .A2(\adder/norm/_0972_ ),
    .A3(\adder/norm/_1006_ ),
    .A4(\adder/norm/_0875_ ),
    .ZN(\adder/norm/_1007_ ));
 NAND3_X1 \adder/norm/_1912_  (.A1(\adder/norm/_0660_ ),
    .A2(net162),
    .A3(net258),
    .ZN(\adder/norm/_1008_ ));
 NOR2_X2 \adder/norm/_1913_  (.A1(\adder/norm/_1008_ ),
    .A2(\adder/norm/_0681_ ),
    .ZN(\adder/norm/_1009_ ));
 NAND3_X1 \adder/norm/_1914_  (.A1(\adder/norm/_1009_ ),
    .A2(\adder/norm/_0694_ ),
    .A3(\adder/norm/_0642_ ),
    .ZN(\adder/norm/_1010_ ));
 OAI21_X1 \adder/norm/_1915_  (.A(\adder/norm/_0892_ ),
    .B1(\adder/norm/_1010_ ),
    .B2(\adder/norm/_0888_ ),
    .ZN(\adder/norm/_1011_ ));
 INV_X1 \adder/norm/_1916_  (.A(\adder/norm/_0650_ ),
    .ZN(\adder/norm/_1012_ ));
 XNOR2_X2 \adder/norm/_1917_  (.A(\adder/norm/_0874_ ),
    .B(\adder/norm/_1012_ ),
    .ZN(\adder/norm/_1013_ ));
 AND2_X1 \adder/norm/_1918_  (.A1(\adder/norm/_1011_ ),
    .A2(\adder/norm/_1013_ ),
    .ZN(\adder/norm/_1014_ ));
 NAND2_X1 \adder/norm/_1919_  (.A1(\adder/norm/_1007_ ),
    .A2(\adder/norm/_1014_ ),
    .ZN(\adder/norm/_1015_ ));
 NOR2_X1 \adder/norm/_1920_  (.A1(\adder/norm/_0896_ ),
    .A2(\adder/norm/_1015_ ),
    .ZN(\adder/norm/_1016_ ));
 NAND2_X1 \adder/norm/_1921_  (.A1(\adder/norm/_0901_ ),
    .A2(\adder/norm/_0681_ ),
    .ZN(\adder/norm/_1017_ ));
 NAND2_X1 \adder/norm/_1922_  (.A1(\adder/norm/_0923_ ),
    .A2(net81),
    .ZN(\adder/norm/_1018_ ));
 TAPCELL_X1 PHY_59 ();
 NAND3_X1 \adder/norm/_1924_  (.A1(\adder/norm/_1017_ ),
    .A2(\adder/norm/_1018_ ),
    .A3(net243),
    .ZN(\adder/norm/_1020_ ));
 NAND3_X1 \adder/norm/_1925_  (.A1(\adder/norm/_0925_ ),
    .A2(\adder/norm/_0926_ ),
    .A3(\adder/norm/_0681_ ),
    .ZN(\adder/norm/_1021_ ));
 NAND3_X1 \adder/norm/_1926_  (.A1(\adder/norm/_0932_ ),
    .A2(net81),
    .A3(\adder/norm/_0933_ ),
    .ZN(\adder/norm/_1022_ ));
 NAND3_X1 \adder/norm/_1927_  (.A1(\adder/norm/_1021_ ),
    .A2(\adder/norm/_1022_ ),
    .A3(\adder/norm/_0694_ ),
    .ZN(\adder/norm/_1023_ ));
 NAND3_X1 \adder/norm/_1928_  (.A1(\adder/norm/_1020_ ),
    .A2(\adder/norm/_1023_ ),
    .A3(net250),
    .ZN(\adder/norm/_1024_ ));
 NAND3_X1 \adder/norm/_1929_  (.A1(\adder/norm/_0909_ ),
    .A2(\adder/norm/_0910_ ),
    .A3(\adder/norm/_0681_ ),
    .ZN(\adder/norm/_1025_ ));
 NAND3_X1 \adder/norm/_1930_  (.A1(\adder/norm/_0903_ ),
    .A2(net81),
    .A3(\adder/norm/_0904_ ),
    .ZN(\adder/norm/_1026_ ));
 NAND3_X1 \adder/norm/_1931_  (.A1(\adder/norm/_1025_ ),
    .A2(\adder/norm/_1026_ ),
    .A3(\adder/norm/_0694_ ),
    .ZN(\adder/norm/_1027_ ));
 NAND3_X1 \adder/norm/_1932_  (.A1(\adder/norm/_0965_ ),
    .A2(\adder/norm/_0966_ ),
    .A3(\adder/norm/_0681_ ),
    .ZN(\adder/norm/_1028_ ));
 NAND3_X1 \adder/norm/_1933_  (.A1(\adder/norm/_0912_ ),
    .A2(\adder/norm/_0913_ ),
    .A3(net81),
    .ZN(\adder/norm/_1029_ ));
 NAND3_X1 \adder/norm/_1934_  (.A1(\adder/norm/_1028_ ),
    .A2(\adder/norm/_1029_ ),
    .A3(net246),
    .ZN(\adder/norm/_1030_ ));
 NAND3_X1 \adder/norm/_1935_  (.A1(\adder/norm/_1027_ ),
    .A2(\adder/norm/_1030_ ),
    .A3(\adder/norm/_0747_ ),
    .ZN(\adder/norm/_1031_ ));
 NAND2_X1 \adder/norm/_1936_  (.A1(\adder/norm/_1024_ ),
    .A2(\adder/norm/_1031_ ),
    .ZN(\adder/norm/_1032_ ));
 NAND2_X1 \adder/norm/_1937_  (.A1(\adder/norm/_1032_ ),
    .A2(\adder/norm/_0761_ ),
    .ZN(\adder/norm/_1033_ ));
 NAND2_X1 \adder/norm/_1938_  (.A1(\adder/norm/_0940_ ),
    .A2(\adder/norm/_0681_ ),
    .ZN(\adder/norm/_1034_ ));
 NAND3_X1 \adder/norm/_1939_  (.A1(\adder/norm/_0946_ ),
    .A2(net81),
    .A3(\adder/norm/_0947_ ),
    .ZN(\adder/norm/_1035_ ));
 NAND3_X1 \adder/norm/_1940_  (.A1(\adder/norm/_1034_ ),
    .A2(\adder/norm/_1035_ ),
    .A3(\adder/norm/_0694_ ),
    .ZN(\adder/norm/_1036_ ));
 NAND3_X1 \adder/norm/_1941_  (.A1(\adder/norm/_0942_ ),
    .A2(net81),
    .A3(\adder/norm/_0943_ ),
    .ZN(\adder/norm/_1037_ ));
 NAND2_X1 \adder/norm/_1942_  (.A1(\adder/norm/_1008_ ),
    .A2(\adder/norm/_0681_ ),
    .ZN(\adder/norm/_1038_ ));
 NAND3_X1 \adder/norm/_1943_  (.A1(\adder/norm/_1037_ ),
    .A2(net246),
    .A3(\adder/norm/_1038_ ),
    .ZN(\adder/norm/_1039_ ));
 NAND3_X1 \adder/norm/_1944_  (.A1(\adder/norm/_1036_ ),
    .A2(\adder/norm/_1039_ ),
    .A3(\adder/norm/_0747_ ),
    .ZN(\adder/norm/_1040_ ));
 NAND3_X1 \adder/norm/_1945_  (.A1(\adder/norm/_0949_ ),
    .A2(\adder/norm/_0681_ ),
    .A3(\adder/norm/_0950_ ),
    .ZN(\adder/norm/_1041_ ));
 NAND3_X1 \adder/norm/_1946_  (.A1(\adder/norm/_0957_ ),
    .A2(\adder/norm/_0958_ ),
    .A3(net81),
    .ZN(\adder/norm/_1042_ ));
 NAND3_X1 \adder/norm/_1947_  (.A1(\adder/norm/_1041_ ),
    .A2(\adder/norm/_1042_ ),
    .A3(net243),
    .ZN(\adder/norm/_1043_ ));
 NAND3_X1 \adder/norm/_1948_  (.A1(\adder/norm/_0954_ ),
    .A2(\adder/norm/_0681_ ),
    .A3(\adder/norm/_0955_ ),
    .ZN(\adder/norm/_1044_ ));
 NAND3_X1 \adder/norm/_1949_  (.A1(\adder/norm/_0962_ ),
    .A2(\adder/norm/_0963_ ),
    .A3(net81),
    .ZN(\adder/norm/_1045_ ));
 NAND3_X1 \adder/norm/_1950_  (.A1(\adder/norm/_1044_ ),
    .A2(\adder/norm/_1045_ ),
    .A3(\adder/norm/_0694_ ),
    .ZN(\adder/norm/_1046_ ));
 NAND3_X1 \adder/norm/_1951_  (.A1(\adder/norm/_1043_ ),
    .A2(\adder/norm/_1046_ ),
    .A3(net250),
    .ZN(\adder/norm/_1047_ ));
 NAND2_X1 \adder/norm/_1952_  (.A1(\adder/norm/_1040_ ),
    .A2(\adder/norm/_1047_ ),
    .ZN(\adder/norm/_1048_ ));
 NAND2_X1 \adder/norm/_1953_  (.A1(\adder/norm/_1048_ ),
    .A2(\adder/norm/_0820_ ),
    .ZN(\adder/norm/_1049_ ));
 NAND2_X1 \adder/norm/_1954_  (.A1(\adder/norm/_1033_ ),
    .A2(\adder/norm/_1049_ ),
    .ZN(\adder/norm/_1050_ ));
 NAND3_X1 \adder/norm/_1955_  (.A1(\adder/norm/_0929_ ),
    .A2(\adder/norm/_0930_ ),
    .A3(\adder/norm/_0681_ ),
    .ZN(\adder/norm/_1051_ ));
 NAND3_X1 \adder/norm/_1956_  (.A1(\adder/norm/_0973_ ),
    .A2(net82),
    .A3(\adder/norm/_0974_ ),
    .ZN(\adder/norm/_1052_ ));
 NAND3_X1 \adder/norm/_1957_  (.A1(\adder/norm/_1051_ ),
    .A2(\adder/norm/_1052_ ),
    .A3(net243),
    .ZN(\adder/norm/_1053_ ));
 NAND3_X1 \adder/norm/_1958_  (.A1(\adder/norm/_0976_ ),
    .A2(\adder/norm/_0681_ ),
    .A3(\adder/norm/_0977_ ),
    .ZN(\adder/norm/_1054_ ));
 NAND3_X1 \adder/norm/_1959_  (.A1(\adder/norm/_0983_ ),
    .A2(\adder/norm/_0984_ ),
    .A3(\adder/norm/_0680_ ),
    .ZN(\adder/norm/_1055_ ));
 NAND3_X1 \adder/norm/_1960_  (.A1(\adder/norm/_1054_ ),
    .A2(\adder/norm/_1055_ ),
    .A3(\adder/norm/_0694_ ),
    .ZN(\adder/norm/_1056_ ));
 NAND3_X1 \adder/norm/_1961_  (.A1(\adder/norm/_1053_ ),
    .A2(\adder/norm/_1056_ ),
    .A3(\adder/norm/_0747_ ),
    .ZN(\adder/norm/_1057_ ));
 NAND3_X1 \adder/norm/_1962_  (.A1(\adder/norm/_0980_ ),
    .A2(\adder/norm/_0681_ ),
    .A3(\adder/norm/_0981_ ),
    .ZN(\adder/norm/_1058_ ));
 NAND3_X1 \adder/norm/_1963_  (.A1(\adder/norm/_0993_ ),
    .A2(\adder/norm/_0994_ ),
    .A3(\adder/norm/_0680_ ),
    .ZN(\adder/norm/_1059_ ));
 NAND3_X1 \adder/norm/_1964_  (.A1(\adder/norm/_1058_ ),
    .A2(\adder/norm/_1059_ ),
    .A3(net243),
    .ZN(\adder/norm/_1060_ ));
 NAND3_X1 \adder/norm/_1965_  (.A1(\adder/norm/_0990_ ),
    .A2(\adder/norm/_0681_ ),
    .A3(\adder/norm/_0991_ ),
    .ZN(\adder/norm/_1061_ ));
 NAND3_X1 \adder/norm/_1966_  (.A1(\adder/norm/_0997_ ),
    .A2(\adder/norm/_0998_ ),
    .A3(\adder/norm/_0680_ ),
    .ZN(\adder/norm/_1062_ ));
 NAND3_X1 \adder/norm/_1967_  (.A1(\adder/norm/_1061_ ),
    .A2(\adder/norm/_1062_ ),
    .A3(\adder/norm/_0694_ ),
    .ZN(\adder/norm/_1063_ ));
 NAND3_X1 \adder/norm/_1968_  (.A1(\adder/norm/_1060_ ),
    .A2(\adder/norm/_1063_ ),
    .A3(net250),
    .ZN(\adder/norm/_1064_ ));
 NAND2_X1 \adder/norm/_1969_  (.A1(\adder/norm/_1057_ ),
    .A2(\adder/norm/_1064_ ),
    .ZN(\adder/norm/_1065_ ));
 NAND2_X1 \adder/norm/_1970_  (.A1(\adder/norm/_1065_ ),
    .A2(\adder/norm/_0870_ ),
    .ZN(\adder/norm/_1066_ ));
 NOR2_X2 \adder/norm/_1971_  (.A1(\adder/norm/_0877_ ),
    .A2(\adder/norm/_0892_ ),
    .ZN(\adder/norm/_1067_ ));
 INV_X2 \adder/norm/_1972_  (.A(\adder/norm/_1067_ ),
    .ZN(\adder/norm/_1068_ ));
 TAPCELL_X1 PHY_58 ();
 NOR2_X1 \adder/norm/_1974_  (.A1(\adder/norm/_1000_ ),
    .A2(\adder/norm/_0680_ ),
    .ZN(\adder/norm/_1070_ ));
 NAND3_X1 \adder/norm/_1975_  (.A1(\adder/norm/_1070_ ),
    .A2(net241),
    .A3(\adder/norm/_0642_ ),
    .ZN(\adder/norm/_1071_ ));
 AOI21_X1 \adder/norm/_1976_  (.A(\adder/norm/_1068_ ),
    .B1(\adder/norm/_1071_ ),
    .B2(\adder/norm/_0889_ ),
    .ZN(\adder/norm/_1072_ ));
 NAND2_X1 \adder/norm/_1977_  (.A1(\adder/norm/_1066_ ),
    .A2(\adder/norm/_1072_ ),
    .ZN(\adder/norm/_1073_ ));
 NOR2_X1 \adder/norm/_1978_  (.A1(\adder/norm/_1050_ ),
    .A2(\adder/norm/_1073_ ),
    .ZN(\adder/norm/_1074_ ));
 NAND2_X1 \adder/norm/_1979_  (.A1(\adder/norm/_0788_ ),
    .A2(\adder/norm/_0681_ ),
    .ZN(\adder/norm/_1075_ ));
 NAND3_X1 \adder/norm/_1980_  (.A1(\adder/norm/_0803_ ),
    .A2(net81),
    .A3(\adder/norm/_0806_ ),
    .ZN(\adder/norm/_1076_ ));
 NAND2_X1 \adder/norm/_1981_  (.A1(\adder/norm/_1075_ ),
    .A2(\adder/norm/_1076_ ),
    .ZN(\adder/norm/_1077_ ));
 NAND2_X1 \adder/norm/_1982_  (.A1(\adder/norm/_1077_ ),
    .A2(net240),
    .ZN(\adder/norm/_1078_ ));
 NAND2_X1 \adder/norm/_1983_  (.A1(\adder/norm/_0801_ ),
    .A2(\adder/norm/_0681_ ),
    .ZN(\adder/norm/_1079_ ));
 NAND3_X1 \adder/norm/_1984_  (.A1(\adder/norm/_0815_ ),
    .A2(net81),
    .A3(\adder/norm/_0816_ ),
    .ZN(\adder/norm/_1080_ ));
 NAND2_X1 \adder/norm/_1985_  (.A1(\adder/norm/_1079_ ),
    .A2(\adder/norm/_1080_ ),
    .ZN(\adder/norm/_1081_ ));
 NAND2_X1 \adder/norm/_1986_  (.A1(\adder/norm/_1081_ ),
    .A2(\adder/norm/_0694_ ),
    .ZN(\adder/norm/_1082_ ));
 NAND3_X1 \adder/norm/_1987_  (.A1(\adder/norm/_1078_ ),
    .A2(\adder/norm/_1082_ ),
    .A3(\adder/norm/_0717_ ),
    .ZN(\adder/norm/_1083_ ));
 NAND2_X1 \adder/norm/_1988_  (.A1(\adder/norm/_0779_ ),
    .A2(\adder/norm/_0681_ ),
    .ZN(\adder/norm/_1084_ ));
 NAND3_X1 \adder/norm/_1989_  (.A1(\adder/norm/_0790_ ),
    .A2(\adder/norm/_0792_ ),
    .A3(net81),
    .ZN(\adder/norm/_1085_ ));
 NAND2_X1 \adder/norm/_1990_  (.A1(\adder/norm/_1084_ ),
    .A2(\adder/norm/_1085_ ),
    .ZN(\adder/norm/_1086_ ));
 NAND2_X1 \adder/norm/_1991_  (.A1(\adder/norm/_1086_ ),
    .A2(\adder/norm/_0694_ ),
    .ZN(\adder/norm/_1087_ ));
 NAND3_X1 \adder/norm/_1992_  (.A1(\adder/norm/_0768_ ),
    .A2(\adder/norm/_0771_ ),
    .A3(net81),
    .ZN(\adder/norm/_1088_ ));
 NAND3_X1 \adder/norm/_1993_  (.A1(\adder/norm/_0879_ ),
    .A2(\adder/norm/_0681_ ),
    .A3(\adder/norm/_0882_ ),
    .ZN(\adder/norm/_1089_ ));
 NAND3_X1 \adder/norm/_1994_  (.A1(\adder/norm/_1088_ ),
    .A2(\adder/norm/_1089_ ),
    .A3(net240),
    .ZN(\adder/norm/_1090_ ));
 NAND3_X1 \adder/norm/_1995_  (.A1(\adder/norm/_1087_ ),
    .A2(\adder/norm/_1090_ ),
    .A3(\adder/norm/_0747_ ),
    .ZN(\adder/norm/_1091_ ));
 NAND3_X1 \adder/norm/_1996_  (.A1(\adder/norm/_1083_ ),
    .A2(\adder/norm/_1091_ ),
    .A3(\adder/norm/_0758_ ),
    .ZN(\adder/norm/_1092_ ));
 NAND2_X1 \adder/norm/_1997_  (.A1(\adder/norm/_0727_ ),
    .A2(\adder/norm/_0681_ ),
    .ZN(\adder/norm/_1093_ ));
 NAND3_X1 \adder/norm/_1998_  (.A1(\adder/norm/_0737_ ),
    .A2(net82),
    .A3(\adder/norm/_0738_ ),
    .ZN(\adder/norm/_1094_ ));
 NAND2_X1 \adder/norm/_1999_  (.A1(\adder/norm/_1093_ ),
    .A2(\adder/norm/_1094_ ),
    .ZN(\adder/norm/_1095_ ));
 NAND2_X1 \adder/norm/_2000_  (.A1(\adder/norm/_1095_ ),
    .A2(\adder/norm/_0694_ ),
    .ZN(\adder/norm/_1096_ ));
 TAPCELL_X1 PHY_57 ();
 INV_X1 \adder/norm/_2002_  (.A(net163),
    .ZN(\adder/norm/_1098_ ));
 OAI21_X1 \adder/norm/_2003_  (.A(\adder/norm/_0673_ ),
    .B1(net247),
    .B2(\adder/norm/_1098_ ),
    .ZN(\adder/norm/_1099_ ));
 INV_X1 \adder/norm/_2004_  (.A(net164),
    .ZN(\adder/norm/_1100_ ));
 OAI21_X1 \adder/norm/_2005_  (.A(net84),
    .B1(net247),
    .B2(\adder/norm/_1100_ ),
    .ZN(\adder/norm/_1101_ ));
 NAND3_X1 \adder/norm/_2006_  (.A1(\adder/norm/_1099_ ),
    .A2(\adder/norm/_1101_ ),
    .A3(net82),
    .ZN(\adder/norm/_1102_ ));
 NAND3_X1 \adder/norm/_2007_  (.A1(\adder/norm/_0810_ ),
    .A2(\adder/norm/_0681_ ),
    .A3(\adder/norm/_0812_ ),
    .ZN(\adder/norm/_1103_ ));
 NAND3_X1 \adder/norm/_2008_  (.A1(\adder/norm/_1102_ ),
    .A2(\adder/norm/_1103_ ),
    .A3(net241),
    .ZN(\adder/norm/_1104_ ));
 NAND3_X1 \adder/norm/_2009_  (.A1(\adder/norm/_1096_ ),
    .A2(\adder/norm/_1104_ ),
    .A3(\adder/norm/_0747_ ),
    .ZN(\adder/norm/_1105_ ));
 NAND3_X1 \adder/norm/_2010_  (.A1(\adder/norm/_0672_ ),
    .A2(\adder/norm/_0677_ ),
    .A3(net82),
    .ZN(\adder/norm/_1106_ ));
 NAND3_X1 \adder/norm/_2011_  (.A1(\adder/norm/_0699_ ),
    .A2(\adder/norm/_0702_ ),
    .A3(\adder/norm/_0681_ ),
    .ZN(\adder/norm/_1107_ ));
 NAND3_X1 \adder/norm/_2012_  (.A1(\adder/norm/_1106_ ),
    .A2(\adder/norm/_1107_ ),
    .A3(\adder/norm/_0694_ ),
    .ZN(\adder/norm/_1108_ ));
 NAND3_X1 \adder/norm/_2013_  (.A1(\adder/norm/_0740_ ),
    .A2(\adder/norm/_0681_ ),
    .A3(\adder/norm/_0741_ ),
    .ZN(\adder/norm/_1109_ ));
 NAND3_X1 \adder/norm/_2014_  (.A1(\adder/norm/_0709_ ),
    .A2(\adder/norm/_0710_ ),
    .A3(net82),
    .ZN(\adder/norm/_1110_ ));
 NAND2_X1 \adder/norm/_2015_  (.A1(\adder/norm/_1109_ ),
    .A2(\adder/norm/_1110_ ),
    .ZN(\adder/norm/_1111_ ));
 NAND2_X1 \adder/norm/_2016_  (.A1(\adder/norm/_1111_ ),
    .A2(net240),
    .ZN(\adder/norm/_1112_ ));
 NAND3_X1 \adder/norm/_2017_  (.A1(\adder/norm/_1108_ ),
    .A2(\adder/norm/_1112_ ),
    .A3(\adder/norm/_0717_ ),
    .ZN(\adder/norm/_1113_ ));
 NAND3_X1 \adder/norm/_2018_  (.A1(\adder/norm/_1105_ ),
    .A2(\adder/norm/_1113_ ),
    .A3(\adder/norm/_0759_ ),
    .ZN(\adder/norm/_1114_ ));
 NAND2_X1 \adder/norm/_2019_  (.A1(\adder/norm/_1092_ ),
    .A2(\adder/norm/_1114_ ),
    .ZN(\adder/norm/_1115_ ));
 NAND2_X1 \adder/norm/_2020_  (.A1(\adder/norm/_1115_ ),
    .A2(\adder/norm/_0755_ ),
    .ZN(\adder/norm/_1116_ ));
 NAND2_X1 \adder/norm/_2021_  (.A1(\adder/norm/_0828_ ),
    .A2(\adder/norm/_0681_ ),
    .ZN(\adder/norm/_1117_ ));
 NAND3_X1 \adder/norm/_2022_  (.A1(\adder/norm/_0855_ ),
    .A2(net82),
    .A3(\adder/norm/_0857_ ),
    .ZN(\adder/norm/_1118_ ));
 NAND3_X1 \adder/norm/_2023_  (.A1(\adder/norm/_1117_ ),
    .A2(\adder/norm/_1118_ ),
    .A3(net243),
    .ZN(\adder/norm/_1119_ ));
 NAND3_X1 \adder/norm/_2024_  (.A1(\adder/norm/_0852_ ),
    .A2(\adder/norm/_0853_ ),
    .A3(\adder/norm/_0681_ ),
    .ZN(\adder/norm/_1120_ ));
 NAND3_X1 \adder/norm/_2025_  (.A1(\adder/norm/_0861_ ),
    .A2(net82),
    .A3(\adder/norm/_0863_ ),
    .ZN(\adder/norm/_1121_ ));
 NAND3_X1 \adder/norm/_2026_  (.A1(\adder/norm/_1120_ ),
    .A2(\adder/norm/_1121_ ),
    .A3(\adder/norm/_0694_ ),
    .ZN(\adder/norm/_1122_ ));
 NAND3_X1 \adder/norm/_2027_  (.A1(\adder/norm/_1119_ ),
    .A2(\adder/norm/_1122_ ),
    .A3(net250),
    .ZN(\adder/norm/_1123_ ));
 NAND3_X1 \adder/norm/_2028_  (.A1(\adder/norm/_0688_ ),
    .A2(\adder/norm/_0691_ ),
    .A3(\adder/norm/_0681_ ),
    .ZN(\adder/norm/_1124_ ));
 NAND3_X1 \adder/norm/_2029_  (.A1(\adder/norm/_0839_ ),
    .A2(net82),
    .A3(\adder/norm/_0840_ ),
    .ZN(\adder/norm/_1125_ ));
 NAND3_X1 \adder/norm/_2030_  (.A1(\adder/norm/_1124_ ),
    .A2(\adder/norm/_1125_ ),
    .A3(net241),
    .ZN(\adder/norm/_1126_ ));
 NAND3_X1 \adder/norm/_2031_  (.A1(\adder/norm/_0845_ ),
    .A2(\adder/norm/_0681_ ),
    .A3(\adder/norm/_0847_ ),
    .ZN(\adder/norm/_1127_ ));
 NAND3_X1 \adder/norm/_2032_  (.A1(\adder/norm/_0834_ ),
    .A2(\adder/norm/_0835_ ),
    .A3(net82),
    .ZN(\adder/norm/_1128_ ));
 NAND3_X1 \adder/norm/_2033_  (.A1(\adder/norm/_1127_ ),
    .A2(\adder/norm/_1128_ ),
    .A3(\adder/norm/_0694_ ),
    .ZN(\adder/norm/_1129_ ));
 NAND3_X1 \adder/norm/_2034_  (.A1(\adder/norm/_1126_ ),
    .A2(\adder/norm/_1129_ ),
    .A3(\adder/norm/_0747_ ),
    .ZN(\adder/norm/_1130_ ));
 NAND3_X1 \adder/norm/_2035_  (.A1(\adder/norm/_1123_ ),
    .A2(\adder/norm/_1130_ ),
    .A3(\adder/norm/_0758_ ),
    .ZN(\adder/norm/_1131_ ));
 AOI21_X1 \adder/norm/_2036_  (.A(\adder/norm/_1068_ ),
    .B1(\adder/norm/_1131_ ),
    .B2(\adder/norm/_0754_ ),
    .ZN(\adder/norm/_1132_ ));
 NAND3_X1 \adder/norm/_2037_  (.A1(\adder/norm/_1074_ ),
    .A2(\adder/norm/_1116_ ),
    .A3(\adder/norm/_1132_ ),
    .ZN(\adder/norm/_1133_ ));
 NAND2_X1 \adder/norm/_2038_  (.A1(\adder/norm/_0774_ ),
    .A2(\adder/norm/_0782_ ),
    .ZN(\adder/norm/_1134_ ));
 NAND2_X1 \adder/norm/_2039_  (.A1(\adder/norm/_1134_ ),
    .A2(\adder/norm/_0694_ ),
    .ZN(\adder/norm/_1135_ ));
 NAND2_X1 \adder/norm/_2040_  (.A1(\adder/norm/_0883_ ),
    .A2(net240),
    .ZN(\adder/norm/_1136_ ));
 NAND2_X1 \adder/norm/_2041_  (.A1(\adder/norm/_1135_ ),
    .A2(\adder/norm/_1136_ ),
    .ZN(\adder/norm/_1137_ ));
 NAND2_X1 \adder/norm/_2042_  (.A1(\adder/norm/_1137_ ),
    .A2(\adder/norm/_0747_ ),
    .ZN(\adder/norm/_1138_ ));
 NAND2_X1 \adder/norm/_2043_  (.A1(\adder/norm/_0789_ ),
    .A2(\adder/norm/_0793_ ),
    .ZN(\adder/norm/_1139_ ));
 NAND2_X1 \adder/norm/_2044_  (.A1(\adder/norm/_1139_ ),
    .A2(net240),
    .ZN(\adder/norm/_1140_ ));
 NAND2_X1 \adder/norm/_2045_  (.A1(\adder/norm/_0802_ ),
    .A2(\adder/norm/_0807_ ),
    .ZN(\adder/norm/_1141_ ));
 NAND2_X1 \adder/norm/_2046_  (.A1(\adder/norm/_1141_ ),
    .A2(\adder/norm/_0694_ ),
    .ZN(\adder/norm/_1142_ ));
 NAND2_X1 \adder/norm/_2047_  (.A1(\adder/norm/_1140_ ),
    .A2(\adder/norm/_1142_ ),
    .ZN(\adder/norm/_1143_ ));
 NAND2_X1 \adder/norm/_2048_  (.A1(\adder/norm/_1143_ ),
    .A2(net250),
    .ZN(\adder/norm/_1144_ ));
 NAND2_X1 \adder/norm/_2049_  (.A1(\adder/norm/_1138_ ),
    .A2(\adder/norm/_1144_ ),
    .ZN(\adder/norm/_1145_ ));
 NAND2_X1 \adder/norm/_2050_  (.A1(\adder/norm/_1145_ ),
    .A2(\adder/norm/_0820_ ),
    .ZN(\adder/norm/_1146_ ));
 NAND2_X1 \adder/norm/_2051_  (.A1(\adder/norm/_0705_ ),
    .A2(\adder/norm/_0712_ ),
    .ZN(\adder/norm/_1147_ ));
 NAND2_X1 \adder/norm/_2052_  (.A1(\adder/norm/_1147_ ),
    .A2(\adder/norm/_0694_ ),
    .ZN(\adder/norm/_1148_ ));
 NAND2_X1 \adder/norm/_2053_  (.A1(\adder/norm/_0743_ ),
    .A2(net240),
    .ZN(\adder/norm/_1149_ ));
 NAND2_X1 \adder/norm/_2054_  (.A1(\adder/norm/_1148_ ),
    .A2(\adder/norm/_1149_ ),
    .ZN(\adder/norm/_1150_ ));
 NAND2_X1 \adder/norm/_2055_  (.A1(\adder/norm/_1150_ ),
    .A2(net250),
    .ZN(\adder/norm/_1151_ ));
 NAND2_X1 \adder/norm/_2056_  (.A1(\adder/norm/_0733_ ),
    .A2(\adder/norm/_0694_ ),
    .ZN(\adder/norm/_1152_ ));
 NAND2_X1 \adder/norm/_2057_  (.A1(\adder/norm/_0814_ ),
    .A2(\adder/norm/_0817_ ),
    .ZN(\adder/norm/_1153_ ));
 NAND2_X1 \adder/norm/_2058_  (.A1(\adder/norm/_1153_ ),
    .A2(net240),
    .ZN(\adder/norm/_1154_ ));
 NAND2_X1 \adder/norm/_2059_  (.A1(\adder/norm/_1152_ ),
    .A2(\adder/norm/_1154_ ),
    .ZN(\adder/norm/_1155_ ));
 NAND2_X1 \adder/norm/_2060_  (.A1(\adder/norm/_1155_ ),
    .A2(\adder/norm/_0747_ ),
    .ZN(\adder/norm/_1156_ ));
 NAND2_X1 \adder/norm/_2061_  (.A1(\adder/norm/_1151_ ),
    .A2(\adder/norm/_1156_ ),
    .ZN(\adder/norm/_1157_ ));
 NAND2_X1 \adder/norm/_2062_  (.A1(\adder/norm/_1157_ ),
    .A2(\adder/norm/_0761_ ),
    .ZN(\adder/norm/_1158_ ));
 NAND2_X1 \adder/norm/_2063_  (.A1(\adder/norm/_1146_ ),
    .A2(\adder/norm/_1158_ ),
    .ZN(\adder/norm/_1159_ ));
 NAND3_X1 \adder/norm/_2064_  (.A1(\adder/norm/_0684_ ),
    .A2(\adder/norm/_0693_ ),
    .A3(net243),
    .ZN(\adder/norm/_1160_ ));
 NAND3_X1 \adder/norm/_2065_  (.A1(\adder/norm/_0841_ ),
    .A2(\adder/norm/_0848_ ),
    .A3(\adder/norm/_0694_ ),
    .ZN(\adder/norm/_1161_ ));
 NAND3_X1 \adder/norm/_2066_  (.A1(\adder/norm/_1160_ ),
    .A2(\adder/norm/_1161_ ),
    .A3(\adder/norm/_0747_ ),
    .ZN(\adder/norm/_1162_ ));
 NAND3_X1 \adder/norm/_2067_  (.A1(\adder/norm/_0829_ ),
    .A2(\adder/norm/_0836_ ),
    .A3(net243),
    .ZN(\adder/norm/_1163_ ));
 NAND3_X1 \adder/norm/_2068_  (.A1(\adder/norm/_0854_ ),
    .A2(\adder/norm/_0858_ ),
    .A3(\adder/norm/_0694_ ),
    .ZN(\adder/norm/_1164_ ));
 NAND3_X1 \adder/norm/_2069_  (.A1(\adder/norm/_1163_ ),
    .A2(\adder/norm/_1164_ ),
    .A3(net250),
    .ZN(\adder/norm/_1165_ ));
 NAND2_X1 \adder/norm/_2070_  (.A1(\adder/norm/_1162_ ),
    .A2(\adder/norm/_1165_ ),
    .ZN(\adder/norm/_1166_ ));
 NAND2_X1 \adder/norm/_2071_  (.A1(\adder/norm/_1166_ ),
    .A2(\adder/norm/_0870_ ),
    .ZN(\adder/norm/_1167_ ));
 NAND4_X1 \adder/norm/_2072_  (.A1(\adder/norm/_0864_ ),
    .A2(net241),
    .A3(\adder/norm/_0642_ ),
    .A4(\adder/norm/_0681_ ),
    .ZN(\adder/norm/_1168_ ));
 AOI21_X1 \adder/norm/_2073_  (.A(\adder/norm/_1068_ ),
    .B1(\adder/norm/_1168_ ),
    .B2(\adder/norm/_0889_ ),
    .ZN(\adder/norm/_1169_ ));
 NAND2_X1 \adder/norm/_2074_  (.A1(\adder/norm/_1167_ ),
    .A2(\adder/norm/_1169_ ),
    .ZN(\adder/norm/_1170_ ));
 NOR2_X1 \adder/norm/_2075_  (.A1(\adder/norm/_1159_ ),
    .A2(\adder/norm/_1170_ ),
    .ZN(\adder/norm/_1171_ ));
 NAND3_X1 \adder/norm/_2076_  (.A1(\adder/norm/_0902_ ),
    .A2(\adder/norm/_0905_ ),
    .A3(net243),
    .ZN(\adder/norm/_1172_ ));
 NAND3_X1 \adder/norm/_2077_  (.A1(\adder/norm/_0924_ ),
    .A2(\adder/norm/_0927_ ),
    .A3(\adder/norm/_0694_ ),
    .ZN(\adder/norm/_1173_ ));
 NAND3_X1 \adder/norm/_2078_  (.A1(\adder/norm/_1172_ ),
    .A2(\adder/norm/_1173_ ),
    .A3(\adder/norm/_0717_ ),
    .ZN(\adder/norm/_1174_ ));
 NAND2_X1 \adder/norm/_2079_  (.A1(\adder/norm/_0915_ ),
    .A2(\adder/norm/_0694_ ),
    .ZN(\adder/norm/_1175_ ));
 NAND2_X1 \adder/norm/_2080_  (.A1(\adder/norm/_0968_ ),
    .A2(net240),
    .ZN(\adder/norm/_1176_ ));
 NAND2_X1 \adder/norm/_2081_  (.A1(\adder/norm/_1175_ ),
    .A2(\adder/norm/_1176_ ),
    .ZN(\adder/norm/_1177_ ));
 NAND2_X1 \adder/norm/_2082_  (.A1(\adder/norm/_1177_ ),
    .A2(\adder/norm/_0747_ ),
    .ZN(\adder/norm/_1178_ ));
 NAND2_X1 \adder/norm/_2083_  (.A1(\adder/norm/_1174_ ),
    .A2(\adder/norm/_1178_ ),
    .ZN(\adder/norm/_1179_ ));
 NAND2_X1 \adder/norm/_2084_  (.A1(\adder/norm/_1179_ ),
    .A2(\adder/norm/_0761_ ),
    .ZN(\adder/norm/_1180_ ));
 NAND3_X1 \adder/norm/_2085_  (.A1(\adder/norm/_0941_ ),
    .A2(\adder/norm/_0944_ ),
    .A3(\adder/norm/_0694_ ),
    .ZN(\adder/norm/_1181_ ));
 TAPCELL_X1 PHY_56 ();
 NAND2_X1 \adder/norm/_2087_  (.A1(\adder/norm/_1009_ ),
    .A2(net240),
    .ZN(\adder/norm/_1183_ ));
 NAND3_X1 \adder/norm/_2088_  (.A1(\adder/norm/_1181_ ),
    .A2(\adder/norm/_0747_ ),
    .A3(\adder/norm/_1183_ ),
    .ZN(\adder/norm/_1184_ ));
 NAND3_X1 \adder/norm/_2089_  (.A1(\adder/norm/_0948_ ),
    .A2(\adder/norm/_0951_ ),
    .A3(net243),
    .ZN(\adder/norm/_1185_ ));
 NAND3_X1 \adder/norm/_2090_  (.A1(\adder/norm/_0956_ ),
    .A2(\adder/norm/_0959_ ),
    .A3(\adder/norm/_0694_ ),
    .ZN(\adder/norm/_1186_ ));
 NAND3_X1 \adder/norm/_2091_  (.A1(\adder/norm/_1185_ ),
    .A2(\adder/norm/_1186_ ),
    .A3(\adder/norm/_0717_ ),
    .ZN(\adder/norm/_1187_ ));
 NAND2_X1 \adder/norm/_2092_  (.A1(\adder/norm/_1184_ ),
    .A2(\adder/norm/_1187_ ),
    .ZN(\adder/norm/_1188_ ));
 NAND2_X1 \adder/norm/_2093_  (.A1(\adder/norm/_1188_ ),
    .A2(\adder/norm/_0820_ ),
    .ZN(\adder/norm/_1189_ ));
 NAND2_X1 \adder/norm/_2094_  (.A1(\adder/norm/_1180_ ),
    .A2(\adder/norm/_1189_ ),
    .ZN(\adder/norm/_1190_ ));
 NAND2_X1 \adder/norm/_2095_  (.A1(\adder/norm/_0931_ ),
    .A2(\adder/norm/_0934_ ),
    .ZN(\adder/norm/_1191_ ));
 NAND2_X1 \adder/norm/_2096_  (.A1(\adder/norm/_1191_ ),
    .A2(net240),
    .ZN(\adder/norm/_1192_ ));
 NAND2_X1 \adder/norm/_2097_  (.A1(\adder/norm/_0975_ ),
    .A2(\adder/norm/_0978_ ),
    .ZN(\adder/norm/_1193_ ));
 NAND2_X1 \adder/norm/_2098_  (.A1(\adder/norm/_1193_ ),
    .A2(\adder/norm/_0694_ ),
    .ZN(\adder/norm/_1194_ ));
 NAND2_X1 \adder/norm/_2099_  (.A1(\adder/norm/_1192_ ),
    .A2(\adder/norm/_1194_ ),
    .ZN(\adder/norm/_1195_ ));
 NAND2_X1 \adder/norm/_2100_  (.A1(\adder/norm/_1195_ ),
    .A2(\adder/norm/_0747_ ),
    .ZN(\adder/norm/_1196_ ));
 NAND2_X1 \adder/norm/_2101_  (.A1(\adder/norm/_0992_ ),
    .A2(\adder/norm/_0995_ ),
    .ZN(\adder/norm/_1197_ ));
 NAND2_X1 \adder/norm/_2102_  (.A1(\adder/norm/_1197_ ),
    .A2(\adder/norm/_0694_ ),
    .ZN(\adder/norm/_1198_ ));
 NAND2_X1 \adder/norm/_2103_  (.A1(\adder/norm/_0982_ ),
    .A2(\adder/norm/_0985_ ),
    .ZN(\adder/norm/_1199_ ));
 NAND2_X1 \adder/norm/_2104_  (.A1(\adder/norm/_1199_ ),
    .A2(net240),
    .ZN(\adder/norm/_1200_ ));
 NAND2_X1 \adder/norm/_2105_  (.A1(\adder/norm/_1198_ ),
    .A2(\adder/norm/_1200_ ),
    .ZN(\adder/norm/_1201_ ));
 NAND2_X1 \adder/norm/_2106_  (.A1(\adder/norm/_1201_ ),
    .A2(net250),
    .ZN(\adder/norm/_1202_ ));
 NAND2_X1 \adder/norm/_2107_  (.A1(\adder/norm/_1196_ ),
    .A2(\adder/norm/_1202_ ),
    .ZN(\adder/norm/_1203_ ));
 NAND2_X1 \adder/norm/_2108_  (.A1(\adder/norm/_1203_ ),
    .A2(\adder/norm/_0870_ ),
    .ZN(\adder/norm/_1204_ ));
 NAND3_X1 \adder/norm/_2109_  (.A1(\adder/norm/_0999_ ),
    .A2(\adder/norm/_1001_ ),
    .A3(net243),
    .ZN(\adder/norm/_1205_ ));
 OR2_X1 \adder/norm/_2110_  (.A1(\adder/norm/_1205_ ),
    .A2(net250),
    .ZN(\adder/norm/_1206_ ));
 AOI21_X1 \adder/norm/_2111_  (.A(\adder/norm/_1068_ ),
    .B1(\adder/norm/_1206_ ),
    .B2(\adder/norm/_0889_ ),
    .ZN(\adder/norm/_1207_ ));
 NAND2_X1 \adder/norm/_2112_  (.A1(\adder/norm/_1204_ ),
    .A2(\adder/norm/_1207_ ),
    .ZN(\adder/norm/_1208_ ));
 NOR2_X2 \adder/norm/_2113_  (.A1(\adder/norm/_1190_ ),
    .A2(\adder/norm/_1208_ ),
    .ZN(\adder/norm/_1209_ ));
 NAND2_X1 \adder/norm/_2114_  (.A1(\adder/norm/_1171_ ),
    .A2(\adder/norm/_1209_ ),
    .ZN(\adder/norm/_1210_ ));
 NOR2_X2 \adder/norm/_2115_  (.A1(\adder/norm/_1133_ ),
    .A2(\adder/norm/_1210_ ),
    .ZN(\adder/norm/_1211_ ));
 NAND2_X1 \adder/norm/_2116_  (.A1(\adder/norm/_1088_ ),
    .A2(\adder/norm/_1089_ ),
    .ZN(\adder/norm/_1212_ ));
 NAND3_X1 \adder/norm/_2117_  (.A1(\adder/norm/_1212_ ),
    .A2(\adder/norm/_0694_ ),
    .A3(\adder/norm/_0642_ ),
    .ZN(\adder/norm/_1213_ ));
 OAI21_X1 \adder/norm/_2118_  (.A(\adder/norm/_0892_ ),
    .B1(\adder/norm/_1213_ ),
    .B2(\adder/norm/_0888_ ),
    .ZN(\adder/norm/_1214_ ));
 AND2_X1 \adder/norm/_2119_  (.A1(\adder/norm/_1214_ ),
    .A2(\adder/norm/_1013_ ),
    .ZN(\adder/norm/_1215_ ));
 NAND3_X1 \adder/norm/_2120_  (.A1(\adder/norm/_1106_ ),
    .A2(\adder/norm/_1107_ ),
    .A3(net240),
    .ZN(\adder/norm/_1216_ ));
 NAND2_X1 \adder/norm/_2121_  (.A1(\adder/norm/_1124_ ),
    .A2(\adder/norm/_1125_ ),
    .ZN(\adder/norm/_1217_ ));
 NAND2_X1 \adder/norm/_2122_  (.A1(\adder/norm/_1217_ ),
    .A2(\adder/norm/_0694_ ),
    .ZN(\adder/norm/_1218_ ));
 NAND2_X1 \adder/norm/_2123_  (.A1(\adder/norm/_1216_ ),
    .A2(\adder/norm/_1218_ ),
    .ZN(\adder/norm/_1219_ ));
 NAND2_X1 \adder/norm/_2124_  (.A1(\adder/norm/_1219_ ),
    .A2(\adder/norm/_0717_ ),
    .ZN(\adder/norm/_1220_ ));
 NAND3_X1 \adder/norm/_2125_  (.A1(\adder/norm/_1093_ ),
    .A2(\adder/norm/_1094_ ),
    .A3(net246),
    .ZN(\adder/norm/_1221_ ));
 NAND3_X1 \adder/norm/_2126_  (.A1(\adder/norm/_1109_ ),
    .A2(\adder/norm/_1110_ ),
    .A3(\adder/norm/_0694_ ),
    .ZN(\adder/norm/_1222_ ));
 NAND3_X1 \adder/norm/_2127_  (.A1(\adder/norm/_1221_ ),
    .A2(\adder/norm/_1222_ ),
    .A3(\adder/norm/_0747_ ),
    .ZN(\adder/norm/_1223_ ));
 NAND3_X1 \adder/norm/_2128_  (.A1(\adder/norm/_1220_ ),
    .A2(\adder/norm/_1223_ ),
    .A3(\adder/norm/_0761_ ),
    .ZN(\adder/norm/_1224_ ));
 NAND3_X1 \adder/norm/_2129_  (.A1(\adder/norm/_1084_ ),
    .A2(\adder/norm/_1085_ ),
    .A3(net246),
    .ZN(\adder/norm/_1225_ ));
 NAND3_X1 \adder/norm/_2130_  (.A1(\adder/norm/_1075_ ),
    .A2(\adder/norm/_1076_ ),
    .A3(\adder/norm/_0694_ ),
    .ZN(\adder/norm/_1226_ ));
 NAND3_X1 \adder/norm/_2131_  (.A1(\adder/norm/_1225_ ),
    .A2(\adder/norm/_1226_ ),
    .A3(\adder/norm/_0747_ ),
    .ZN(\adder/norm/_1227_ ));
 NAND3_X1 \adder/norm/_2132_  (.A1(\adder/norm/_1079_ ),
    .A2(\adder/norm/_1080_ ),
    .A3(net246),
    .ZN(\adder/norm/_1228_ ));
 NAND2_X1 \adder/norm/_2133_  (.A1(\adder/norm/_0813_ ),
    .A2(\adder/norm/_0681_ ),
    .ZN(\adder/norm/_1229_ ));
 NAND3_X1 \adder/norm/_2134_  (.A1(\adder/norm/_0730_ ),
    .A2(\adder/norm/_0731_ ),
    .A3(net81),
    .ZN(\adder/norm/_1230_ ));
 NAND3_X1 \adder/norm/_2135_  (.A1(\adder/norm/_1229_ ),
    .A2(\adder/norm/_1230_ ),
    .A3(\adder/norm/_0694_ ),
    .ZN(\adder/norm/_1231_ ));
 TAPCELL_X1 PHY_55 ();
 NAND3_X1 \adder/norm/_2137_  (.A1(\adder/norm/_1228_ ),
    .A2(\adder/norm/_1231_ ),
    .A3(\adder/norm/_0717_ ),
    .ZN(\adder/norm/_1233_ ));
 NAND3_X1 \adder/norm/_2138_  (.A1(\adder/norm/_1227_ ),
    .A2(\adder/norm/_1233_ ),
    .A3(\adder/norm/_0820_ ),
    .ZN(\adder/norm/_1234_ ));
 NAND3_X1 \adder/norm/_2139_  (.A1(\adder/norm/_1117_ ),
    .A2(\adder/norm/_1118_ ),
    .A3(\adder/norm/_0694_ ),
    .ZN(\adder/norm/_1235_ ));
 NAND3_X1 \adder/norm/_2140_  (.A1(\adder/norm/_1127_ ),
    .A2(\adder/norm/_1128_ ),
    .A3(net246),
    .ZN(\adder/norm/_1236_ ));
 NAND3_X1 \adder/norm/_2141_  (.A1(\adder/norm/_1235_ ),
    .A2(\adder/norm/_1236_ ),
    .A3(\adder/norm/_0747_ ),
    .ZN(\adder/norm/_1237_ ));
 NAND2_X1 \adder/norm/_2142_  (.A1(\adder/norm/_1120_ ),
    .A2(\adder/norm/_1121_ ),
    .ZN(\adder/norm/_1238_ ));
 INV_X1 \adder/norm/_2143_  (.A(\adder/norm/_1238_ ),
    .ZN(\adder/norm/_1239_ ));
 NAND2_X1 \adder/norm/_2144_  (.A1(\adder/norm/_1239_ ),
    .A2(net243),
    .ZN(\adder/norm/_1240_ ));
 NAND2_X1 \adder/norm/_2145_  (.A1(\adder/norm/_1240_ ),
    .A2(\adder/norm/_0717_ ),
    .ZN(\adder/norm/_1241_ ));
 NAND3_X1 \adder/norm/_2146_  (.A1(\adder/norm/_1237_ ),
    .A2(\adder/norm/_1241_ ),
    .A3(\adder/norm/_0870_ ),
    .ZN(\adder/norm/_1242_ ));
 NAND3_X1 \adder/norm/_2147_  (.A1(\adder/norm/_1224_ ),
    .A2(\adder/norm/_1234_ ),
    .A3(\adder/norm/_1242_ ),
    .ZN(\adder/norm/_1243_ ));
 OAI21_X1 \adder/norm/_2148_  (.A(\adder/norm/_1215_ ),
    .B1(\adder/norm/_1243_ ),
    .B2(\adder/norm/_0892_ ),
    .ZN(\adder/norm/_1244_ ));
 NAND3_X1 \adder/norm/_2149_  (.A1(\adder/norm/_1017_ ),
    .A2(\adder/norm/_1018_ ),
    .A3(\adder/norm/_0694_ ),
    .ZN(\adder/norm/_1245_ ));
 NAND3_X1 \adder/norm/_2150_  (.A1(\adder/norm/_1025_ ),
    .A2(\adder/norm/_1026_ ),
    .A3(net241),
    .ZN(\adder/norm/_1246_ ));
 NAND3_X1 \adder/norm/_2151_  (.A1(\adder/norm/_1245_ ),
    .A2(\adder/norm/_1246_ ),
    .A3(\adder/norm/_0747_ ),
    .ZN(\adder/norm/_1247_ ));
 NAND3_X1 \adder/norm/_2152_  (.A1(\adder/norm/_1021_ ),
    .A2(\adder/norm/_1022_ ),
    .A3(net241),
    .ZN(\adder/norm/_1248_ ));
 NAND3_X1 \adder/norm/_2153_  (.A1(\adder/norm/_1051_ ),
    .A2(\adder/norm/_1052_ ),
    .A3(\adder/norm/_0694_ ),
    .ZN(\adder/norm/_1249_ ));
 NAND3_X1 \adder/norm/_2154_  (.A1(\adder/norm/_1248_ ),
    .A2(\adder/norm/_1249_ ),
    .A3(\adder/norm/_0717_ ),
    .ZN(\adder/norm/_1250_ ));
 NAND3_X1 \adder/norm/_2155_  (.A1(\adder/norm/_1247_ ),
    .A2(\adder/norm/_1250_ ),
    .A3(\adder/norm/_0761_ ),
    .ZN(\adder/norm/_1251_ ));
 NAND3_X1 \adder/norm/_2156_  (.A1(\adder/norm/_1034_ ),
    .A2(\adder/norm/_1035_ ),
    .A3(net241),
    .ZN(\adder/norm/_1252_ ));
 NAND3_X1 \adder/norm/_2157_  (.A1(\adder/norm/_1041_ ),
    .A2(\adder/norm/_1042_ ),
    .A3(\adder/norm/_0694_ ),
    .ZN(\adder/norm/_1253_ ));
 NAND3_X1 \adder/norm/_2158_  (.A1(\adder/norm/_1252_ ),
    .A2(\adder/norm/_1253_ ),
    .A3(\adder/norm/_0747_ ),
    .ZN(\adder/norm/_1254_ ));
 NAND3_X1 \adder/norm/_2159_  (.A1(\adder/norm/_1044_ ),
    .A2(\adder/norm/_1045_ ),
    .A3(net241),
    .ZN(\adder/norm/_1255_ ));
 NAND3_X1 \adder/norm/_2160_  (.A1(\adder/norm/_1028_ ),
    .A2(\adder/norm/_1029_ ),
    .A3(\adder/norm/_0694_ ),
    .ZN(\adder/norm/_1256_ ));
 NAND3_X1 \adder/norm/_2161_  (.A1(\adder/norm/_1255_ ),
    .A2(\adder/norm/_1256_ ),
    .A3(\adder/norm/_0717_ ),
    .ZN(\adder/norm/_1257_ ));
 NAND3_X1 \adder/norm/_2162_  (.A1(\adder/norm/_1254_ ),
    .A2(\adder/norm/_1257_ ),
    .A3(\adder/norm/_0820_ ),
    .ZN(\adder/norm/_1258_ ));
 NAND3_X1 \adder/norm/_2163_  (.A1(\adder/norm/_1054_ ),
    .A2(\adder/norm/_1055_ ),
    .A3(net241),
    .ZN(\adder/norm/_1259_ ));
 NAND3_X1 \adder/norm/_2164_  (.A1(\adder/norm/_1058_ ),
    .A2(\adder/norm/_1059_ ),
    .A3(\adder/norm/_0694_ ),
    .ZN(\adder/norm/_1260_ ));
 NAND3_X1 \adder/norm/_2165_  (.A1(\adder/norm/_1259_ ),
    .A2(\adder/norm/_1260_ ),
    .A3(\adder/norm/_0747_ ),
    .ZN(\adder/norm/_1261_ ));
 NAND3_X1 \adder/norm/_2166_  (.A1(\adder/norm/_1061_ ),
    .A2(\adder/norm/_1062_ ),
    .A3(net241),
    .ZN(\adder/norm/_1262_ ));
 NAND2_X1 \adder/norm/_2167_  (.A1(\adder/norm/_1070_ ),
    .A2(\adder/norm/_0694_ ),
    .ZN(\adder/norm/_1263_ ));
 NAND3_X1 \adder/norm/_2168_  (.A1(\adder/norm/_1262_ ),
    .A2(\adder/norm/_0717_ ),
    .A3(\adder/norm/_1263_ ),
    .ZN(\adder/norm/_1264_ ));
 NAND3_X1 \adder/norm/_2169_  (.A1(\adder/norm/_1261_ ),
    .A2(\adder/norm/_1264_ ),
    .A3(\adder/norm/_0870_ ),
    .ZN(\adder/norm/_1265_ ));
 NAND4_X1 \adder/norm/_2170_  (.A1(\adder/norm/_1251_ ),
    .A2(\adder/norm/_1258_ ),
    .A3(\adder/norm/_1265_ ),
    .A4(\adder/norm/_0875_ ),
    .ZN(\adder/norm/_1266_ ));
 NAND3_X1 \adder/norm/_2171_  (.A1(\adder/norm/_1037_ ),
    .A2(\adder/norm/_0694_ ),
    .A3(\adder/norm/_1038_ ),
    .ZN(\adder/norm/_1267_ ));
 NOR2_X1 \adder/norm/_2172_  (.A1(\adder/norm/_1267_ ),
    .A2(\adder/norm/_0747_ ),
    .ZN(\adder/norm/_1268_ ));
 NAND2_X1 \adder/norm/_2173_  (.A1(\adder/norm/_1268_ ),
    .A2(\adder/norm/_0889_ ),
    .ZN(\adder/norm/_1269_ ));
 AOI21_X1 \adder/norm/_2174_  (.A(\adder/norm/_0877_ ),
    .B1(\adder/norm/_1269_ ),
    .B2(\adder/norm/_0892_ ),
    .ZN(\adder/norm/_1270_ ));
 NAND2_X1 \adder/norm/_2175_  (.A1(\adder/norm/_1266_ ),
    .A2(\adder/norm/_1270_ ),
    .ZN(\adder/norm/_1271_ ));
 NOR2_X1 \adder/norm/_2176_  (.A1(\adder/norm/_1244_ ),
    .A2(\adder/norm/_1271_ ),
    .ZN(\adder/norm/_1272_ ));
 NAND3_X1 \adder/norm/_2177_  (.A1(\adder/norm/_1016_ ),
    .A2(\adder/norm/_1211_ ),
    .A3(\adder/norm/_1272_ ),
    .ZN(\adder/norm/_1273_ ));
 TAPCELL_X1 PHY_54 ();
 NAND3_X1 \adder/norm/_2179_  (.A1(\adder/norm/_1135_ ),
    .A2(\adder/norm/_1136_ ),
    .A3(\adder/norm/_0717_ ),
    .ZN(\adder/norm/_1275_ ));
 AOI21_X1 \adder/norm/_2180_  (.A(\adder/norm/_1068_ ),
    .B1(\adder/norm/_1275_ ),
    .B2(\adder/norm/_0820_ ),
    .ZN(\adder/norm/_1276_ ));
 NAND2_X1 \adder/norm/_2181_  (.A1(\adder/norm/_1150_ ),
    .A2(\adder/norm/_0747_ ),
    .ZN(\adder/norm/_1277_ ));
 NAND3_X1 \adder/norm/_2182_  (.A1(\adder/norm/_1160_ ),
    .A2(\adder/norm/_1161_ ),
    .A3(\adder/norm/_0717_ ),
    .ZN(\adder/norm/_1278_ ));
 NAND2_X1 \adder/norm/_2183_  (.A1(\adder/norm/_1277_ ),
    .A2(\adder/norm/_1278_ ),
    .ZN(\adder/norm/_1279_ ));
 NAND2_X1 \adder/norm/_2184_  (.A1(\adder/norm/_1279_ ),
    .A2(\adder/norm/_0870_ ),
    .ZN(\adder/norm/_1280_ ));
 NAND2_X1 \adder/norm/_2185_  (.A1(\adder/norm/_1276_ ),
    .A2(\adder/norm/_1280_ ),
    .ZN(\adder/norm/_1281_ ));
 NAND2_X1 \adder/norm/_2186_  (.A1(\adder/norm/_1143_ ),
    .A2(\adder/norm/_0747_ ),
    .ZN(\adder/norm/_1282_ ));
 NAND2_X1 \adder/norm/_2187_  (.A1(\adder/norm/_1155_ ),
    .A2(\adder/norm/_0717_ ),
    .ZN(\adder/norm/_1283_ ));
 NAND2_X1 \adder/norm/_2188_  (.A1(\adder/norm/_1282_ ),
    .A2(\adder/norm/_1283_ ),
    .ZN(\adder/norm/_1284_ ));
 NAND2_X1 \adder/norm/_2189_  (.A1(\adder/norm/_1284_ ),
    .A2(\adder/norm/_0761_ ),
    .ZN(\adder/norm/_1285_ ));
 NAND3_X1 \adder/norm/_2190_  (.A1(\adder/norm/_1163_ ),
    .A2(\adder/norm/_1164_ ),
    .A3(\adder/norm/_0747_ ),
    .ZN(\adder/norm/_1286_ ));
 NAND2_X1 \adder/norm/_2191_  (.A1(\adder/norm/_0864_ ),
    .A2(\adder/norm/_0681_ ),
    .ZN(\adder/norm/_1287_ ));
 OAI21_X1 \adder/norm/_2192_  (.A(\adder/norm/_0717_ ),
    .B1(\adder/norm/_1287_ ),
    .B2(\adder/norm/_0694_ ),
    .ZN(\adder/norm/_1288_ ));
 NAND2_X1 \adder/norm/_2193_  (.A1(\adder/norm/_1286_ ),
    .A2(\adder/norm/_1288_ ),
    .ZN(\adder/norm/_1289_ ));
 NAND2_X1 \adder/norm/_2194_  (.A1(\adder/norm/_1289_ ),
    .A2(\adder/norm/_0889_ ),
    .ZN(\adder/norm/_1290_ ));
 NAND2_X1 \adder/norm/_2195_  (.A1(\adder/norm/_1285_ ),
    .A2(\adder/norm/_1290_ ),
    .ZN(\adder/norm/_1291_ ));
 NOR2_X2 \adder/norm/_2196_  (.A1(\adder/norm/_1281_ ),
    .A2(\adder/norm/_1291_ ),
    .ZN(\adder/norm/_1292_ ));
 NAND3_X1 \adder/norm/_2197_  (.A1(\adder/norm/_1172_ ),
    .A2(\adder/norm/_1173_ ),
    .A3(\adder/norm/_0747_ ),
    .ZN(\adder/norm/_1293_ ));
 NAND2_X1 \adder/norm/_2198_  (.A1(\adder/norm/_1195_ ),
    .A2(\adder/norm/_0717_ ),
    .ZN(\adder/norm/_1294_ ));
 NAND2_X1 \adder/norm/_2199_  (.A1(\adder/norm/_1293_ ),
    .A2(\adder/norm/_1294_ ),
    .ZN(\adder/norm/_1295_ ));
 NAND2_X1 \adder/norm/_2200_  (.A1(\adder/norm/_1295_ ),
    .A2(\adder/norm/_0870_ ),
    .ZN(\adder/norm/_1296_ ));
 NAND2_X1 \adder/norm/_2201_  (.A1(\adder/norm/_1181_ ),
    .A2(\adder/norm/_1183_ ),
    .ZN(\adder/norm/_1297_ ));
 NAND2_X1 \adder/norm/_2202_  (.A1(\adder/norm/_1297_ ),
    .A2(\adder/norm/_0717_ ),
    .ZN(\adder/norm/_1298_ ));
 AOI21_X1 \adder/norm/_2203_  (.A(\adder/norm/_1068_ ),
    .B1(\adder/norm/_1298_ ),
    .B2(\adder/norm/_0820_ ),
    .ZN(\adder/norm/_1299_ ));
 NAND2_X1 \adder/norm/_2204_  (.A1(\adder/norm/_1296_ ),
    .A2(\adder/norm/_1299_ ),
    .ZN(\adder/norm/_1300_ ));
 NAND2_X1 \adder/norm/_2205_  (.A1(\adder/norm/_1177_ ),
    .A2(\adder/norm/_0717_ ),
    .ZN(\adder/norm/_1301_ ));
 NAND3_X1 \adder/norm/_2206_  (.A1(\adder/norm/_1185_ ),
    .A2(\adder/norm/_1186_ ),
    .A3(\adder/norm/_0747_ ),
    .ZN(\adder/norm/_1302_ ));
 NAND2_X1 \adder/norm/_2207_  (.A1(\adder/norm/_1301_ ),
    .A2(\adder/norm/_1302_ ),
    .ZN(\adder/norm/_1303_ ));
 NAND2_X1 \adder/norm/_2208_  (.A1(\adder/norm/_1303_ ),
    .A2(\adder/norm/_0761_ ),
    .ZN(\adder/norm/_1304_ ));
 NAND2_X1 \adder/norm/_2209_  (.A1(\adder/norm/_1201_ ),
    .A2(\adder/norm/_0747_ ),
    .ZN(\adder/norm/_1305_ ));
 NAND2_X1 \adder/norm/_2210_  (.A1(\adder/norm/_1205_ ),
    .A2(\adder/norm/_0717_ ),
    .ZN(\adder/norm/_1306_ ));
 NAND2_X1 \adder/norm/_2211_  (.A1(\adder/norm/_1305_ ),
    .A2(\adder/norm/_1306_ ),
    .ZN(\adder/norm/_1307_ ));
 NAND2_X1 \adder/norm/_2212_  (.A1(\adder/norm/_1307_ ),
    .A2(\adder/norm/_0889_ ),
    .ZN(\adder/norm/_1308_ ));
 NAND2_X1 \adder/norm/_2213_  (.A1(\adder/norm/_1304_ ),
    .A2(\adder/norm/_1308_ ),
    .ZN(\adder/norm/_1309_ ));
 NOR2_X2 \adder/norm/_2214_  (.A1(\adder/norm/_1300_ ),
    .A2(\adder/norm/_1309_ ),
    .ZN(\adder/norm/_1310_ ));
 NAND2_X1 \adder/norm/_2215_  (.A1(\adder/norm/_1220_ ),
    .A2(\adder/norm/_1223_ ),
    .ZN(\adder/norm/_1311_ ));
 NAND2_X1 \adder/norm/_2216_  (.A1(\adder/norm/_1311_ ),
    .A2(\adder/norm/_0870_ ),
    .ZN(\adder/norm/_1312_ ));
 AOI21_X1 \adder/norm/_2217_  (.A(\adder/norm/_1068_ ),
    .B1(\adder/norm/_1213_ ),
    .B2(\adder/norm/_0820_ ),
    .ZN(\adder/norm/_1313_ ));
 NAND2_X1 \adder/norm/_2218_  (.A1(\adder/norm/_1312_ ),
    .A2(\adder/norm/_1313_ ),
    .ZN(\adder/norm/_1314_ ));
 NAND2_X1 \adder/norm/_2219_  (.A1(\adder/norm/_1227_ ),
    .A2(\adder/norm/_1233_ ),
    .ZN(\adder/norm/_1315_ ));
 NAND2_X1 \adder/norm/_2220_  (.A1(\adder/norm/_1315_ ),
    .A2(\adder/norm/_0761_ ),
    .ZN(\adder/norm/_1316_ ));
 NAND2_X1 \adder/norm/_2221_  (.A1(\adder/norm/_1237_ ),
    .A2(\adder/norm/_1241_ ),
    .ZN(\adder/norm/_1317_ ));
 NAND2_X1 \adder/norm/_2222_  (.A1(\adder/norm/_1317_ ),
    .A2(\adder/norm/_0889_ ),
    .ZN(\adder/norm/_1318_ ));
 NAND2_X1 \adder/norm/_2223_  (.A1(\adder/norm/_1316_ ),
    .A2(\adder/norm/_1318_ ),
    .ZN(\adder/norm/_1319_ ));
 NOR2_X4 \adder/norm/_2224_  (.A1(\adder/norm/_1314_ ),
    .A2(\adder/norm/_1319_ ),
    .ZN(\adder/norm/_1320_ ));
 NAND3_X2 \adder/norm/_2225_  (.A1(\adder/norm/_1292_ ),
    .A2(\adder/norm/_1310_ ),
    .A3(\adder/norm/_1320_ ),
    .ZN(\adder/norm/_1321_ ));
 NAND2_X1 \adder/norm/_2226_  (.A1(\adder/norm/_1078_ ),
    .A2(\adder/norm/_1082_ ),
    .ZN(\adder/norm/_1322_ ));
 NAND2_X1 \adder/norm/_2227_  (.A1(\adder/norm/_1322_ ),
    .A2(\adder/norm/_0747_ ),
    .ZN(\adder/norm/_1323_ ));
 NAND2_X1 \adder/norm/_2228_  (.A1(\adder/norm/_1096_ ),
    .A2(\adder/norm/_1104_ ),
    .ZN(\adder/norm/_1324_ ));
 NAND2_X1 \adder/norm/_2229_  (.A1(\adder/norm/_1324_ ),
    .A2(\adder/norm/_0717_ ),
    .ZN(\adder/norm/_1325_ ));
 NAND2_X1 \adder/norm/_2230_  (.A1(\adder/norm/_1323_ ),
    .A2(\adder/norm/_1325_ ),
    .ZN(\adder/norm/_1326_ ));
 NAND2_X1 \adder/norm/_2231_  (.A1(\adder/norm/_1326_ ),
    .A2(\adder/norm/_0761_ ),
    .ZN(\adder/norm/_1327_ ));
 NAND2_X1 \adder/norm/_2232_  (.A1(\adder/norm/_1108_ ),
    .A2(\adder/norm/_1112_ ),
    .ZN(\adder/norm/_1328_ ));
 NAND2_X1 \adder/norm/_2233_  (.A1(\adder/norm/_1328_ ),
    .A2(\adder/norm/_0747_ ),
    .ZN(\adder/norm/_1329_ ));
 NAND3_X1 \adder/norm/_2234_  (.A1(\adder/norm/_1126_ ),
    .A2(\adder/norm/_1129_ ),
    .A3(\adder/norm/_0717_ ),
    .ZN(\adder/norm/_1330_ ));
 AND2_X1 \adder/norm/_2235_  (.A1(\adder/norm/_1329_ ),
    .A2(\adder/norm/_1330_ ),
    .ZN(\adder/norm/_1331_ ));
 OAI21_X1 \adder/norm/_2236_  (.A(\adder/norm/_1327_ ),
    .B1(\adder/norm/_0869_ ),
    .B2(\adder/norm/_1331_ ),
    .ZN(\adder/norm/_1332_ ));
 NAND2_X1 \adder/norm/_2237_  (.A1(\adder/norm/_1119_ ),
    .A2(\adder/norm/_1122_ ),
    .ZN(\adder/norm/_1333_ ));
 INV_X1 \adder/norm/_2238_  (.A(\adder/norm/_1333_ ),
    .ZN(\adder/norm/_1334_ ));
 OAI21_X1 \adder/norm/_2239_  (.A(\adder/norm/_0889_ ),
    .B1(\adder/norm/_1334_ ),
    .B2(net250),
    .ZN(\adder/norm/_1335_ ));
 NAND3_X1 \adder/norm/_2240_  (.A1(\adder/norm/_1087_ ),
    .A2(\adder/norm/_0717_ ),
    .A3(\adder/norm/_1090_ ),
    .ZN(\adder/norm/_1336_ ));
 NAND2_X1 \adder/norm/_2241_  (.A1(\adder/norm/_1336_ ),
    .A2(\adder/norm/_0820_ ),
    .ZN(\adder/norm/_1337_ ));
 NAND3_X1 \adder/norm/_2242_  (.A1(\adder/norm/_1335_ ),
    .A2(\adder/norm/_1067_ ),
    .A3(\adder/norm/_1337_ ),
    .ZN(\adder/norm/_1338_ ));
 NOR2_X2 \adder/norm/_2243_  (.A1(\adder/norm/_1332_ ),
    .A2(\adder/norm/_1338_ ),
    .ZN(\adder/norm/_1339_ ));
 NAND2_X1 \adder/norm/_2244_  (.A1(\adder/norm/_1036_ ),
    .A2(\adder/norm/_1039_ ),
    .ZN(\adder/norm/_1340_ ));
 NAND2_X1 \adder/norm/_2245_  (.A1(\adder/norm/_1340_ ),
    .A2(\adder/norm/_0717_ ),
    .ZN(\adder/norm/_1341_ ));
 AOI21_X1 \adder/norm/_2246_  (.A(\adder/norm/_1068_ ),
    .B1(\adder/norm/_1341_ ),
    .B2(\adder/norm/_0820_ ),
    .ZN(\adder/norm/_1342_ ));
 NAND3_X1 \adder/norm/_2247_  (.A1(\adder/norm/_1020_ ),
    .A2(\adder/norm/_1023_ ),
    .A3(\adder/norm/_0747_ ),
    .ZN(\adder/norm/_1343_ ));
 NAND3_X1 \adder/norm/_2248_  (.A1(\adder/norm/_1053_ ),
    .A2(\adder/norm/_1056_ ),
    .A3(\adder/norm/_0717_ ),
    .ZN(\adder/norm/_1344_ ));
 AND2_X1 \adder/norm/_2249_  (.A1(\adder/norm/_1343_ ),
    .A2(\adder/norm/_1344_ ),
    .ZN(\adder/norm/_1345_ ));
 OAI21_X1 \adder/norm/_2250_  (.A(\adder/norm/_1342_ ),
    .B1(\adder/norm/_0869_ ),
    .B2(\adder/norm/_1345_ ),
    .ZN(\adder/norm/_1346_ ));
 NAND3_X1 \adder/norm/_2251_  (.A1(\adder/norm/_1027_ ),
    .A2(\adder/norm/_1030_ ),
    .A3(\adder/norm/_0717_ ),
    .ZN(\adder/norm/_1347_ ));
 NAND3_X1 \adder/norm/_2252_  (.A1(\adder/norm/_1043_ ),
    .A2(\adder/norm/_1046_ ),
    .A3(\adder/norm/_0747_ ),
    .ZN(\adder/norm/_1348_ ));
 NAND2_X1 \adder/norm/_2253_  (.A1(\adder/norm/_1347_ ),
    .A2(\adder/norm/_1348_ ),
    .ZN(\adder/norm/_1349_ ));
 NAND2_X1 \adder/norm/_2254_  (.A1(\adder/norm/_1349_ ),
    .A2(\adder/norm/_0761_ ),
    .ZN(\adder/norm/_1350_ ));
 NAND3_X1 \adder/norm/_2255_  (.A1(\adder/norm/_1060_ ),
    .A2(\adder/norm/_1063_ ),
    .A3(\adder/norm/_0747_ ),
    .ZN(\adder/norm/_1351_ ));
 INV_X1 \adder/norm/_2256_  (.A(\adder/norm/_1070_ ),
    .ZN(\adder/norm/_1352_ ));
 OAI21_X1 \adder/norm/_2257_  (.A(\adder/norm/_0717_ ),
    .B1(\adder/norm/_1352_ ),
    .B2(\adder/norm/_0694_ ),
    .ZN(\adder/norm/_1353_ ));
 AND2_X1 \adder/norm/_2258_  (.A1(\adder/norm/_1351_ ),
    .A2(\adder/norm/_1353_ ),
    .ZN(\adder/norm/_1354_ ));
 OAI21_X1 \adder/norm/_2259_  (.A(\adder/norm/_1350_ ),
    .B1(\adder/norm/_1354_ ),
    .B2(\adder/norm/_0888_ ),
    .ZN(\adder/norm/_1355_ ));
 NOR2_X2 \adder/norm/_2260_  (.A1(\adder/norm/_1346_ ),
    .A2(\adder/norm/_1355_ ),
    .ZN(\adder/norm/_1356_ ));
 NAND2_X1 \adder/norm/_2261_  (.A1(\adder/norm/_1339_ ),
    .A2(\adder/norm/_1356_ ),
    .ZN(\adder/norm/_1357_ ));
 NOR2_X4 \adder/norm/_2262_  (.A1(\adder/norm/_1357_ ),
    .A2(\adder/norm/_1321_ ),
    .ZN(\adder/norm/_1358_ ));
 NAND2_X1 \adder/norm/_2263_  (.A1(\adder/norm/_0854_ ),
    .A2(\adder/norm/_0858_ ),
    .ZN(\adder/norm/_1359_ ));
 NAND2_X1 \adder/norm/_2264_  (.A1(\adder/norm/_1359_ ),
    .A2(net240),
    .ZN(\adder/norm/_1360_ ));
 NAND2_X1 \adder/norm/_2265_  (.A1(\adder/norm/_1287_ ),
    .A2(\adder/norm/_0694_ ),
    .ZN(\adder/norm/_1361_ ));
 NAND3_X1 \adder/norm/_2266_  (.A1(\adder/norm/_1360_ ),
    .A2(\adder/norm/_0747_ ),
    .A3(\adder/norm/_1361_ ),
    .ZN(\adder/norm/_1362_ ));
 AOI21_X1 \adder/norm/_2267_  (.A(\adder/norm/_1068_ ),
    .B1(\adder/norm/_1362_ ),
    .B2(\adder/norm/_0889_ ),
    .ZN(\adder/norm/_1363_ ));
 NAND2_X1 \adder/norm/_2268_  (.A1(\adder/norm/_0714_ ),
    .A2(\adder/norm/_0747_ ),
    .ZN(\adder/norm/_1364_ ));
 NAND3_X1 \adder/norm/_2269_  (.A1(\adder/norm/_0838_ ),
    .A2(\adder/norm/_0850_ ),
    .A3(\adder/norm/_0717_ ),
    .ZN(\adder/norm/_1365_ ));
 NAND2_X1 \adder/norm/_2270_  (.A1(\adder/norm/_1364_ ),
    .A2(\adder/norm/_1365_ ),
    .ZN(\adder/norm/_1366_ ));
 INV_X1 \adder/norm/_2271_  (.A(\adder/norm/_1366_ ),
    .ZN(\adder/norm/_1367_ ));
 OAI21_X1 \adder/norm/_2272_  (.A(\adder/norm/_1363_ ),
    .B1(\adder/norm/_1367_ ),
    .B2(\adder/norm/_0869_ ),
    .ZN(\adder/norm/_1368_ ));
 NAND2_X1 \adder/norm/_2273_  (.A1(\adder/norm/_0746_ ),
    .A2(net250),
    .ZN(\adder/norm/_1369_ ));
 NAND3_X1 \adder/norm/_2274_  (.A1(\adder/norm/_0808_ ),
    .A2(\adder/norm/_0818_ ),
    .A3(\adder/norm/_0747_ ),
    .ZN(\adder/norm/_1370_ ));
 AOI21_X1 \adder/norm/_2275_  (.A(\adder/norm/_0760_ ),
    .B1(\adder/norm/_1369_ ),
    .B2(\adder/norm/_1370_ ),
    .ZN(\adder/norm/_1371_ ));
 INV_X2 \adder/norm/_2276_  (.A(\adder/norm/_0820_ ),
    .ZN(\adder/norm/_1372_ ));
 NAND3_X1 \adder/norm/_2277_  (.A1(\adder/norm/_0783_ ),
    .A2(\adder/norm/_0795_ ),
    .A3(\adder/norm/_0717_ ),
    .ZN(\adder/norm/_1373_ ));
 NAND2_X1 \adder/norm/_2278_  (.A1(\adder/norm/_0886_ ),
    .A2(\adder/norm/_0747_ ),
    .ZN(\adder/norm/_1374_ ));
 AOI21_X1 \adder/norm/_2279_  (.A(\adder/norm/_1372_ ),
    .B1(\adder/norm/_1373_ ),
    .B2(\adder/norm/_1374_ ),
    .ZN(\adder/norm/_1375_ ));
 OR2_X1 \adder/norm/_2280_  (.A1(\adder/norm/_1371_ ),
    .A2(\adder/norm/_1375_ ),
    .ZN(\adder/norm/_1376_ ));
 NOR2_X4 \adder/norm/_2281_  (.A1(\adder/norm/_1376_ ),
    .A2(\adder/norm/_1368_ ),
    .ZN(\adder/norm/_1377_ ));
 NAND2_X1 \adder/norm/_2282_  (.A1(\adder/norm/_0917_ ),
    .A2(\adder/norm/_0717_ ),
    .ZN(\adder/norm/_1378_ ));
 NAND2_X1 \adder/norm/_2283_  (.A1(\adder/norm/_0970_ ),
    .A2(\adder/norm/_0747_ ),
    .ZN(\adder/norm/_1379_ ));
 AOI21_X1 \adder/norm/_2284_  (.A(\adder/norm/_0760_ ),
    .B1(\adder/norm/_1378_ ),
    .B2(\adder/norm/_1379_ ),
    .ZN(\adder/norm/_1380_ ));
 NAND3_X1 \adder/norm/_2285_  (.A1(\adder/norm/_0945_ ),
    .A2(\adder/norm/_0952_ ),
    .A3(\adder/norm/_0717_ ),
    .ZN(\adder/norm/_1381_ ));
 INV_X1 \adder/norm/_2286_  (.A(\adder/norm/_1009_ ),
    .ZN(\adder/norm/_1382_ ));
 OAI21_X1 \adder/norm/_2287_  (.A(\adder/norm/_0747_ ),
    .B1(\adder/norm/_1382_ ),
    .B2(net240),
    .ZN(\adder/norm/_1383_ ));
 AOI21_X1 \adder/norm/_2288_  (.A(\adder/norm/_1372_ ),
    .B1(\adder/norm/_1381_ ),
    .B2(\adder/norm/_1383_ ),
    .ZN(\adder/norm/_1384_ ));
 OR2_X1 \adder/norm/_2289_  (.A1(\adder/norm/_1380_ ),
    .A2(\adder/norm/_1384_ ),
    .ZN(\adder/norm/_1385_ ));
 NAND2_X1 \adder/norm/_2290_  (.A1(\adder/norm/_0996_ ),
    .A2(\adder/norm/_1002_ ),
    .ZN(\adder/norm/_1386_ ));
 NAND2_X1 \adder/norm/_2291_  (.A1(\adder/norm/_1386_ ),
    .A2(\adder/norm/_0747_ ),
    .ZN(\adder/norm/_1387_ ));
 AOI21_X1 \adder/norm/_2292_  (.A(\adder/norm/_1068_ ),
    .B1(\adder/norm/_1387_ ),
    .B2(\adder/norm/_0889_ ),
    .ZN(\adder/norm/_1388_ ));
 NAND3_X1 \adder/norm/_2293_  (.A1(\adder/norm/_0928_ ),
    .A2(\adder/norm/_0935_ ),
    .A3(\adder/norm/_0747_ ),
    .ZN(\adder/norm/_1389_ ));
 NAND3_X1 \adder/norm/_2294_  (.A1(\adder/norm/_0979_ ),
    .A2(\adder/norm/_0986_ ),
    .A3(\adder/norm/_0717_ ),
    .ZN(\adder/norm/_1390_ ));
 NAND2_X1 \adder/norm/_2295_  (.A1(\adder/norm/_1389_ ),
    .A2(\adder/norm/_1390_ ),
    .ZN(\adder/norm/_1391_ ));
 INV_X1 \adder/norm/_2296_  (.A(\adder/norm/_1391_ ),
    .ZN(\adder/norm/_1392_ ));
 OAI21_X1 \adder/norm/_2297_  (.A(\adder/norm/_1388_ ),
    .B1(\adder/norm/_1392_ ),
    .B2(\adder/norm/_0869_ ),
    .ZN(\adder/norm/_1393_ ));
 NOR2_X4 \adder/norm/_2298_  (.A1(\adder/norm/_1385_ ),
    .A2(\adder/norm/_1393_ ),
    .ZN(\adder/norm/_1394_ ));
 NAND2_X1 \adder/norm/_2299_  (.A1(\adder/norm/_1377_ ),
    .A2(\adder/norm/_1394_ ),
    .ZN(\adder/norm/_1395_ ));
 NAND3_X1 \adder/norm/_2300_  (.A1(\adder/norm/_1228_ ),
    .A2(\adder/norm/_1231_ ),
    .A3(\adder/norm/_0747_ ),
    .ZN(\adder/norm/_1396_ ));
 NAND3_X1 \adder/norm/_2301_  (.A1(\adder/norm/_1221_ ),
    .A2(\adder/norm/_1222_ ),
    .A3(\adder/norm/_0717_ ),
    .ZN(\adder/norm/_1397_ ));
 AOI21_X1 \adder/norm/_2302_  (.A(\adder/norm/_0760_ ),
    .B1(\adder/norm/_1396_ ),
    .B2(\adder/norm/_1397_ ),
    .ZN(\adder/norm/_1398_ ));
 NAND3_X1 \adder/norm/_2303_  (.A1(\adder/norm/_1225_ ),
    .A2(\adder/norm/_1226_ ),
    .A3(\adder/norm/_0717_ ),
    .ZN(\adder/norm/_1399_ ));
 INV_X1 \adder/norm/_2304_  (.A(\adder/norm/_1212_ ),
    .ZN(\adder/norm/_1400_ ));
 OAI21_X1 \adder/norm/_2305_  (.A(\adder/norm/_0747_ ),
    .B1(\adder/norm/_1400_ ),
    .B2(net240),
    .ZN(\adder/norm/_1401_ ));
 AOI21_X1 \adder/norm/_2306_  (.A(\adder/norm/_1372_ ),
    .B1(\adder/norm/_1399_ ),
    .B2(\adder/norm/_1401_ ),
    .ZN(\adder/norm/_1402_ ));
 OR2_X1 \adder/norm/_2307_  (.A1(\adder/norm/_1398_ ),
    .A2(\adder/norm/_1402_ ),
    .ZN(\adder/norm/_1403_ ));
 NAND2_X1 \adder/norm/_2308_  (.A1(\adder/norm/_1219_ ),
    .A2(\adder/norm/_0747_ ),
    .ZN(\adder/norm/_1404_ ));
 NAND3_X1 \adder/norm/_2309_  (.A1(\adder/norm/_1235_ ),
    .A2(\adder/norm/_1236_ ),
    .A3(\adder/norm/_0717_ ),
    .ZN(\adder/norm/_1405_ ));
 NAND2_X1 \adder/norm/_2310_  (.A1(\adder/norm/_1404_ ),
    .A2(\adder/norm/_1405_ ),
    .ZN(\adder/norm/_1406_ ));
 NAND2_X1 \adder/norm/_2311_  (.A1(\adder/norm/_1406_ ),
    .A2(\adder/norm/_0870_ ),
    .ZN(\adder/norm/_1407_ ));
 OAI21_X1 \adder/norm/_2312_  (.A(\adder/norm/_0889_ ),
    .B1(\adder/norm/_1240_ ),
    .B2(net250),
    .ZN(\adder/norm/_1408_ ));
 NAND3_X1 \adder/norm/_2313_  (.A1(\adder/norm/_1407_ ),
    .A2(\adder/norm/_1067_ ),
    .A3(\adder/norm/_1408_ ),
    .ZN(\adder/norm/_1409_ ));
 NOR2_X2 \adder/norm/_2314_  (.A1(\adder/norm/_1403_ ),
    .A2(\adder/norm/_1409_ ),
    .ZN(\adder/norm/_1410_ ));
 NAND3_X1 \adder/norm/_2315_  (.A1(\adder/norm/_1245_ ),
    .A2(\adder/norm/_1246_ ),
    .A3(\adder/norm/_0717_ ),
    .ZN(\adder/norm/_1411_ ));
 NAND3_X1 \adder/norm/_2316_  (.A1(\adder/norm/_1255_ ),
    .A2(\adder/norm/_1256_ ),
    .A3(\adder/norm/_0747_ ),
    .ZN(\adder/norm/_1412_ ));
 AOI21_X1 \adder/norm/_2317_  (.A(\adder/norm/_0760_ ),
    .B1(\adder/norm/_1411_ ),
    .B2(\adder/norm/_1412_ ),
    .ZN(\adder/norm/_1413_ ));
 NAND3_X1 \adder/norm/_2318_  (.A1(\adder/norm/_1252_ ),
    .A2(\adder/norm/_1253_ ),
    .A3(\adder/norm/_0717_ ),
    .ZN(\adder/norm/_1414_ ));
 NAND2_X1 \adder/norm/_2319_  (.A1(\adder/norm/_1267_ ),
    .A2(\adder/norm/_0747_ ),
    .ZN(\adder/norm/_1415_ ));
 AOI21_X1 \adder/norm/_2320_  (.A(\adder/norm/_1372_ ),
    .B1(\adder/norm/_1414_ ),
    .B2(\adder/norm/_1415_ ),
    .ZN(\adder/norm/_1416_ ));
 OR2_X1 \adder/norm/_2321_  (.A1(\adder/norm/_1413_ ),
    .A2(\adder/norm/_1416_ ),
    .ZN(\adder/norm/_1417_ ));
 NAND2_X1 \adder/norm/_2322_  (.A1(\adder/norm/_1262_ ),
    .A2(\adder/norm/_1263_ ),
    .ZN(\adder/norm/_1418_ ));
 NAND2_X1 \adder/norm/_2323_  (.A1(\adder/norm/_1418_ ),
    .A2(\adder/norm/_0747_ ),
    .ZN(\adder/norm/_1419_ ));
 AOI21_X1 \adder/norm/_2324_  (.A(\adder/norm/_1068_ ),
    .B1(\adder/norm/_1419_ ),
    .B2(\adder/norm/_0889_ ),
    .ZN(\adder/norm/_1420_ ));
 NAND3_X1 \adder/norm/_2325_  (.A1(\adder/norm/_1248_ ),
    .A2(\adder/norm/_1249_ ),
    .A3(\adder/norm/_0747_ ),
    .ZN(\adder/norm/_1421_ ));
 NAND3_X1 \adder/norm/_2326_  (.A1(\adder/norm/_1259_ ),
    .A2(\adder/norm/_1260_ ),
    .A3(\adder/norm/_0717_ ),
    .ZN(\adder/norm/_1422_ ));
 NAND2_X1 \adder/norm/_2327_  (.A1(\adder/norm/_1421_ ),
    .A2(\adder/norm/_1422_ ),
    .ZN(\adder/norm/_1423_ ));
 INV_X1 \adder/norm/_2328_  (.A(\adder/norm/_1423_ ),
    .ZN(\adder/norm/_1424_ ));
 OAI21_X1 \adder/norm/_2329_  (.A(\adder/norm/_1420_ ),
    .B1(\adder/norm/_1424_ ),
    .B2(\adder/norm/_0869_ ),
    .ZN(\adder/norm/_1425_ ));
 NOR2_X2 \adder/norm/_2330_  (.A1(\adder/norm/_1417_ ),
    .A2(\adder/norm/_1425_ ),
    .ZN(\adder/norm/_1426_ ));
 NAND2_X1 \adder/norm/_2331_  (.A1(\adder/norm/_1410_ ),
    .A2(\adder/norm/_1426_ ),
    .ZN(\adder/norm/_1427_ ));
 NOR2_X2 \adder/norm/_2332_  (.A1(\adder/norm/_1395_ ),
    .A2(\adder/norm/_1427_ ),
    .ZN(\adder/norm/_1428_ ));
 NAND2_X2 \adder/norm/_2333_  (.A1(\adder/norm/_1358_ ),
    .A2(\adder/norm/_1428_ ),
    .ZN(\adder/norm/_1429_ ));
 NOR2_X4 \adder/norm/_2334_  (.A1(\adder/norm/_1429_ ),
    .A2(\adder/norm/_1273_ ),
    .ZN(\adder/norm/_1430_ ));
 INV_X1 \adder/norm/_2335_  (.A(\adder/mant_prenorm_d[46] ),
    .ZN(\adder/norm/_1431_ ));
 OAI21_X2 \adder/norm/_2336_  (.A(\adder/norm/_0021_ ),
    .B1(\adder/norm/_0666_ ),
    .B2(\adder/norm/_1431_ ),
    .ZN(\adder/norm/_1432_ ));
 XNOR2_X2 \adder/norm/_2337_  (.A(\adder/norm/_1432_ ),
    .B(\adder/norm/Mant_leadingOne_D[0] ),
    .ZN(\adder/norm/_1433_ ));
 NAND3_X1 \adder/norm/_2338_  (.A1(\adder/norm/_1404_ ),
    .A2(\adder/norm/_1405_ ),
    .A3(\adder/norm/_0761_ ),
    .ZN(\adder/norm/_1434_ ));
 NAND3_X1 \adder/norm/_2339_  (.A1(\adder/norm/_1396_ ),
    .A2(\adder/norm/_1397_ ),
    .A3(\adder/norm/_0820_ ),
    .ZN(\adder/norm/_1435_ ));
 NAND4_X1 \adder/norm/_2340_  (.A1(\adder/norm/_1239_ ),
    .A2(net241),
    .A3(\adder/norm/_0747_ ),
    .A4(\adder/norm/_0870_ ),
    .ZN(\adder/norm/_1436_ ));
 NAND3_X1 \adder/norm/_2341_  (.A1(\adder/norm/_1434_ ),
    .A2(\adder/norm/_1435_ ),
    .A3(\adder/norm/_1436_ ),
    .ZN(\adder/norm/_1437_ ));
 NAND2_X1 \adder/norm/_2342_  (.A1(\adder/norm/_1437_ ),
    .A2(\adder/norm/_0875_ ),
    .ZN(\adder/norm/_1438_ ));
 NAND4_X1 \adder/norm/_2343_  (.A1(\adder/norm/_1399_ ),
    .A2(\adder/norm/_1401_ ),
    .A3(\adder/norm/_0892_ ),
    .A4(\adder/norm/_0889_ ),
    .ZN(\adder/norm/_1439_ ));
 NAND2_X1 \adder/norm/_2344_  (.A1(\adder/norm/_1438_ ),
    .A2(\adder/norm/_1439_ ),
    .ZN(\adder/norm/_1440_ ));
 NAND2_X1 \adder/norm/_2345_  (.A1(\adder/norm/_1440_ ),
    .A2(\adder/norm/_1013_ ),
    .ZN(\adder/norm/_1441_ ));
 NAND3_X1 \adder/norm/_2346_  (.A1(\adder/norm/_1414_ ),
    .A2(\adder/norm/_0889_ ),
    .A3(\adder/norm/_1415_ ),
    .ZN(\adder/norm/_1442_ ));
 AOI21_X1 \adder/norm/_2347_  (.A(\adder/norm/_0877_ ),
    .B1(\adder/norm/_1442_ ),
    .B2(\adder/norm/_0892_ ),
    .ZN(\adder/norm/_1443_ ));
 NAND2_X1 \adder/norm/_2348_  (.A1(\adder/norm/_1424_ ),
    .A2(\adder/norm/_0761_ ),
    .ZN(\adder/norm/_1444_ ));
 TAPCELL_X1 PHY_53 ();
 NAND3_X1 \adder/norm/_2350_  (.A1(\adder/norm/_1418_ ),
    .A2(\adder/norm/_0747_ ),
    .A3(\adder/norm/_0870_ ),
    .ZN(\adder/norm/_1446_ ));
 NAND3_X1 \adder/norm/_2351_  (.A1(\adder/norm/_1411_ ),
    .A2(\adder/norm/_1412_ ),
    .A3(\adder/norm/_0820_ ),
    .ZN(\adder/norm/_1447_ ));
 NAND3_X1 \adder/norm/_2352_  (.A1(\adder/norm/_1444_ ),
    .A2(\adder/norm/_1446_ ),
    .A3(\adder/norm/_1447_ ),
    .ZN(\adder/norm/_1448_ ));
 OAI21_X1 \adder/norm/_2353_  (.A(\adder/norm/_1443_ ),
    .B1(\adder/norm/_1448_ ),
    .B2(\adder/norm/_0892_ ),
    .ZN(\adder/norm/_1449_ ));
 NOR2_X1 \adder/norm/_2354_  (.A1(\adder/norm/_1441_ ),
    .A2(\adder/norm/_1449_ ),
    .ZN(\adder/norm/_1450_ ));
 NAND3_X1 \adder/norm/_2355_  (.A1(\adder/norm/_1373_ ),
    .A2(\adder/norm/_0889_ ),
    .A3(\adder/norm/_1374_ ),
    .ZN(\adder/norm/_1451_ ));
 AOI21_X1 \adder/norm/_2356_  (.A(\adder/norm/_0877_ ),
    .B1(\adder/norm/_1451_ ),
    .B2(\adder/norm/_0892_ ),
    .ZN(\adder/norm/_1452_ ));
 NAND3_X1 \adder/norm/_2357_  (.A1(\adder/norm/_1364_ ),
    .A2(\adder/norm/_1365_ ),
    .A3(\adder/norm/_0761_ ),
    .ZN(\adder/norm/_1453_ ));
 OR2_X1 \adder/norm/_2358_  (.A1(\adder/norm/_1362_ ),
    .A2(\adder/norm/_0869_ ),
    .ZN(\adder/norm/_1454_ ));
 NAND3_X1 \adder/norm/_2359_  (.A1(\adder/norm/_1369_ ),
    .A2(\adder/norm/_1370_ ),
    .A3(\adder/norm/_0820_ ),
    .ZN(\adder/norm/_1455_ ));
 NAND3_X1 \adder/norm/_2360_  (.A1(\adder/norm/_1453_ ),
    .A2(\adder/norm/_1454_ ),
    .A3(\adder/norm/_1455_ ),
    .ZN(\adder/norm/_1456_ ));
 OAI21_X1 \adder/norm/_2361_  (.A(\adder/norm/_1452_ ),
    .B1(\adder/norm/_1456_ ),
    .B2(\adder/norm/_0892_ ),
    .ZN(\adder/norm/_1457_ ));
 NAND3_X1 \adder/norm/_2362_  (.A1(\adder/norm/_1381_ ),
    .A2(\adder/norm/_0889_ ),
    .A3(\adder/norm/_1383_ ),
    .ZN(\adder/norm/_1458_ ));
 AOI21_X1 \adder/norm/_2363_  (.A(\adder/norm/_0877_ ),
    .B1(\adder/norm/_1458_ ),
    .B2(\adder/norm/_0892_ ),
    .ZN(\adder/norm/_1459_ ));
 NAND2_X1 \adder/norm/_2364_  (.A1(\adder/norm/_1392_ ),
    .A2(\adder/norm/_0761_ ),
    .ZN(\adder/norm/_1460_ ));
 NAND3_X1 \adder/norm/_2365_  (.A1(\adder/norm/_1378_ ),
    .A2(\adder/norm/_1379_ ),
    .A3(\adder/norm/_0820_ ),
    .ZN(\adder/norm/_1461_ ));
 NAND3_X1 \adder/norm/_2366_  (.A1(\adder/norm/_1386_ ),
    .A2(\adder/norm/_0747_ ),
    .A3(\adder/norm/_0870_ ),
    .ZN(\adder/norm/_1462_ ));
 NAND3_X1 \adder/norm/_2367_  (.A1(\adder/norm/_1460_ ),
    .A2(\adder/norm/_1461_ ),
    .A3(\adder/norm/_1462_ ),
    .ZN(\adder/norm/_1463_ ));
 OAI21_X2 \adder/norm/_2368_  (.A(\adder/norm/_1459_ ),
    .B1(\adder/norm/_1463_ ),
    .B2(\adder/norm/_0892_ ),
    .ZN(\adder/norm/_1465_ ));
 NOR2_X1 \adder/norm/_2369_  (.A1(\adder/norm/_1457_ ),
    .A2(\adder/norm/_1465_ ),
    .ZN(\adder/norm/_1466_ ));
 NAND2_X1 \adder/norm/_2370_  (.A1(\adder/norm/_1450_ ),
    .A2(\adder/norm/_1466_ ),
    .ZN(\adder/norm/_1467_ ));
 OAI21_X1 \adder/norm/_2371_  (.A(\adder/norm/_0892_ ),
    .B1(\adder/norm/_1275_ ),
    .B2(\adder/norm/_0888_ ),
    .ZN(\adder/norm/_1468_ ));
 NAND2_X1 \adder/norm/_2372_  (.A1(\adder/norm/_1468_ ),
    .A2(\adder/norm/_1013_ ),
    .ZN(\adder/norm/_1469_ ));
 INV_X1 \adder/norm/_2373_  (.A(\adder/norm/_1469_ ),
    .ZN(\adder/norm/_1470_ ));
 NAND3_X1 \adder/norm/_2374_  (.A1(\adder/norm/_1282_ ),
    .A2(\adder/norm/_1283_ ),
    .A3(\adder/norm/_0820_ ),
    .ZN(\adder/norm/_1471_ ));
 NAND3_X1 \adder/norm/_2375_  (.A1(\adder/norm/_1277_ ),
    .A2(\adder/norm/_1278_ ),
    .A3(\adder/norm/_0761_ ),
    .ZN(\adder/norm/_1472_ ));
 NAND3_X1 \adder/norm/_2376_  (.A1(\adder/norm/_1286_ ),
    .A2(\adder/norm/_0870_ ),
    .A3(\adder/norm/_1288_ ),
    .ZN(\adder/norm/_1473_ ));
 NAND3_X1 \adder/norm/_2377_  (.A1(\adder/norm/_1471_ ),
    .A2(\adder/norm/_1472_ ),
    .A3(\adder/norm/_1473_ ),
    .ZN(\adder/norm/_1474_ ));
 OAI21_X1 \adder/norm/_2378_  (.A(\adder/norm/_1470_ ),
    .B1(\adder/norm/_1474_ ),
    .B2(\adder/norm/_0892_ ),
    .ZN(\adder/norm/_0000_ ));
 OAI21_X1 \adder/norm/_2379_  (.A(\adder/norm/_0892_ ),
    .B1(\adder/norm/_1298_ ),
    .B2(\adder/norm/_0888_ ),
    .ZN(\adder/norm/_0001_ ));
 NAND2_X1 \adder/norm/_2380_  (.A1(\adder/norm/_0001_ ),
    .A2(\adder/norm/_1013_ ),
    .ZN(\adder/norm/_0002_ ));
 INV_X1 \adder/norm/_2381_  (.A(\adder/norm/_0002_ ),
    .ZN(\adder/norm/_0003_ ));
 NAND3_X1 \adder/norm/_2382_  (.A1(\adder/norm/_1293_ ),
    .A2(\adder/norm/_1294_ ),
    .A3(\adder/norm/_0761_ ),
    .ZN(\adder/norm/_0004_ ));
 NAND3_X1 \adder/norm/_2383_  (.A1(\adder/norm/_1301_ ),
    .A2(\adder/norm/_0820_ ),
    .A3(\adder/norm/_1302_ ),
    .ZN(\adder/norm/_0005_ ));
 NAND3_X1 \adder/norm/_2384_  (.A1(\adder/norm/_1305_ ),
    .A2(\adder/norm/_0870_ ),
    .A3(\adder/norm/_1306_ ),
    .ZN(\adder/norm/_0006_ ));
 NAND3_X1 \adder/norm/_2385_  (.A1(\adder/norm/_0004_ ),
    .A2(\adder/norm/_0005_ ),
    .A3(\adder/norm/_0006_ ),
    .ZN(\adder/norm/_0007_ ));
 OAI21_X1 \adder/norm/_2386_  (.A(\adder/norm/_0003_ ),
    .B1(\adder/norm/_0007_ ),
    .B2(\adder/norm/_0892_ ),
    .ZN(\adder/norm/_0008_ ));
 NOR2_X1 \adder/norm/_2387_  (.A1(\adder/norm/_0000_ ),
    .A2(\adder/norm/_0008_ ),
    .ZN(\adder/norm/_0009_ ));
 OAI21_X1 \adder/norm/_2388_  (.A(\adder/norm/_0892_ ),
    .B1(\adder/norm/_1336_ ),
    .B2(\adder/norm/_0888_ ),
    .ZN(\adder/norm/_0011_ ));
 NAND2_X1 \adder/norm/_2389_  (.A1(\adder/norm/_0011_ ),
    .A2(\adder/norm/_1013_ ),
    .ZN(\adder/norm/_0012_ ));
 INV_X1 \adder/norm/_2390_  (.A(\adder/norm/_0012_ ),
    .ZN(\adder/norm/_0013_ ));
 NAND3_X1 \adder/norm/_2391_  (.A1(\adder/norm/_1323_ ),
    .A2(\adder/norm/_1325_ ),
    .A3(\adder/norm/_0820_ ),
    .ZN(\adder/norm/_0014_ ));
 NAND3_X1 \adder/norm/_2392_  (.A1(\adder/norm/_1329_ ),
    .A2(\adder/norm/_1330_ ),
    .A3(\adder/norm/_0761_ ),
    .ZN(\adder/norm/_0015_ ));
 NAND3_X1 \adder/norm/_2393_  (.A1(\adder/norm/_1333_ ),
    .A2(\adder/norm/_0747_ ),
    .A3(\adder/norm/_0870_ ),
    .ZN(\adder/norm/_0016_ ));
 NAND3_X1 \adder/norm/_2394_  (.A1(\adder/norm/_0014_ ),
    .A2(\adder/norm/_0015_ ),
    .A3(\adder/norm/_0016_ ),
    .ZN(\adder/norm/_0017_ ));
 OAI21_X1 \adder/norm/_2395_  (.A(\adder/norm/_0013_ ),
    .B1(\adder/norm/_0017_ ),
    .B2(\adder/norm/_0892_ ),
    .ZN(\adder/norm/_0018_ ));
 OAI21_X1 \adder/norm/_2396_  (.A(\adder/norm/_0892_ ),
    .B1(\adder/norm/_1341_ ),
    .B2(\adder/norm/_0888_ ),
    .ZN(\adder/norm/_0019_ ));
 NAND2_X1 \adder/norm/_2397_  (.A1(\adder/norm/_0019_ ),
    .A2(\adder/norm/_1013_ ),
    .ZN(\adder/norm/_0020_ ));
 INV_X1 \adder/norm/_2398_  (.A(\adder/norm/_0020_ ),
    .ZN(\adder/norm/_0022_ ));
 NAND3_X1 \adder/norm/_2399_  (.A1(\adder/norm/_1343_ ),
    .A2(\adder/norm/_1344_ ),
    .A3(\adder/norm/_0761_ ),
    .ZN(\adder/norm/_0023_ ));
 NAND3_X1 \adder/norm/_2400_  (.A1(\adder/norm/_1347_ ),
    .A2(\adder/norm/_1348_ ),
    .A3(\adder/norm/_0820_ ),
    .ZN(\adder/norm/_0024_ ));
 NAND3_X1 \adder/norm/_2401_  (.A1(\adder/norm/_1351_ ),
    .A2(\adder/norm/_0870_ ),
    .A3(\adder/norm/_1353_ ),
    .ZN(\adder/norm/_0025_ ));
 NAND3_X1 \adder/norm/_2402_  (.A1(\adder/norm/_0023_ ),
    .A2(\adder/norm/_0024_ ),
    .A3(\adder/norm/_0025_ ),
    .ZN(\adder/norm/_0026_ ));
 OAI21_X1 \adder/norm/_2403_  (.A(\adder/norm/_0022_ ),
    .B1(\adder/norm/_0026_ ),
    .B2(\adder/norm/_0892_ ),
    .ZN(\adder/norm/_0027_ ));
 NOR2_X1 \adder/norm/_2404_  (.A1(\adder/norm/_0018_ ),
    .A2(\adder/norm/_0027_ ),
    .ZN(\adder/norm/_0028_ ));
 NAND2_X1 \adder/norm/_2405_  (.A1(\adder/norm/_0009_ ),
    .A2(\adder/norm/_0028_ ),
    .ZN(\adder/norm/_0029_ ));
 NOR2_X1 \adder/norm/_2406_  (.A1(\adder/norm/_1467_ ),
    .A2(\adder/norm/_0029_ ),
    .ZN(\adder/norm/_0030_ ));
 NAND3_X1 \adder/norm/_2407_  (.A1(\adder/norm/_1430_ ),
    .A2(\adder/norm/_1433_ ),
    .A3(\adder/norm/_0030_ ),
    .ZN(\adder/norm/_0031_ ));
 INV_X1 \adder/norm/_2408_  (.A(\adder/norm/Mant_leadingOne_D[0] ),
    .ZN(\adder/norm/_0033_ ));
 INV_X1 \adder/norm/_2409_  (.A(\adder/norm/_1475_ ),
    .ZN(\adder/norm/_0034_ ));
 OR2_X1 \adder/norm/_2410_  (.A1(\adder/norm/_0034_ ),
    .A2(\adder/norm/_0010_ ),
    .ZN(\adder/norm/_0035_ ));
 NAND3_X1 \adder/norm/_2411_  (.A1(\adder/norm/_1432_ ),
    .A2(\adder/norm/_0033_ ),
    .A3(\adder/norm/_0035_ ),
    .ZN(\adder/norm/_0036_ ));
 INV_X1 \adder/norm/_2412_  (.A(\adder/norm/_0036_ ),
    .ZN(\adder/norm/_0037_ ));
 AOI21_X1 \adder/norm/_2413_  (.A(\adder/norm/_0035_ ),
    .B1(\adder/norm/_1432_ ),
    .B2(\adder/norm/_0033_ ),
    .ZN(\adder/norm/_0038_ ));
 NOR2_X1 \adder/norm/_2414_  (.A1(\adder/norm/_0037_ ),
    .A2(\adder/norm/_0038_ ),
    .ZN(\adder/norm/_0039_ ));
 XNOR2_X1 \adder/norm/_2415_  (.A(\adder/norm/_0031_ ),
    .B(\adder/norm/_0039_ ),
    .ZN(net65));
 NAND4_X1 \adder/norm/_2416_  (.A1(\adder/norm/_1430_ ),
    .A2(\adder/norm/_0030_ ),
    .A3(\adder/norm/_0039_ ),
    .A4(\adder/norm/_1433_ ),
    .ZN(\adder/norm/_0040_ ));
 NAND2_X2 \adder/norm/_2417_  (.A1(\adder/norm/_0040_ ),
    .A2(\adder/norm/_0036_ ),
    .ZN(\adder/norm/_0041_ ));
 XNOR2_X2 \adder/norm/_2418_  (.A(\adder/norm/_0101_ ),
    .B(\adder/norm/_0034_ ),
    .ZN(\adder/norm/_0043_ ));
 XNOR2_X1 \adder/norm/_2419_  (.A(\adder/norm/_0041_ ),
    .B(\adder/norm/_0043_ ),
    .ZN(net66));
 NOR2_X1 \adder/norm/_2420_  (.A1(\adder/norm/_0101_ ),
    .A2(\adder/norm/_0034_ ),
    .ZN(\adder/norm/_0044_ ));
 INV_X1 \adder/norm/_2421_  (.A(\adder/norm/_0043_ ),
    .ZN(\adder/norm/_0045_ ));
 AOI21_X1 \adder/norm/_2422_  (.A(\adder/norm/_0044_ ),
    .B1(\adder/norm/_0041_ ),
    .B2(\adder/norm/_0045_ ),
    .ZN(\adder/norm/_0046_ ));
 XNOR2_X1 \adder/norm/_2423_  (.A(\adder/norm/_0156_ ),
    .B(\adder/norm/_0090_ ),
    .ZN(\adder/norm/_0047_ ));
 INV_X1 \adder/norm/_2424_  (.A(\adder/norm/_0047_ ),
    .ZN(\adder/norm/_0048_ ));
 XNOR2_X1 \adder/norm/_2425_  (.A(\adder/norm/_0046_ ),
    .B(\adder/norm/_0048_ ),
    .ZN(net67));
 NOR2_X1 \adder/norm/_2426_  (.A1(\adder/norm/_0043_ ),
    .A2(\adder/norm/_0047_ ),
    .ZN(\adder/norm/_0049_ ));
 NAND2_X1 \adder/norm/_2427_  (.A1(\adder/norm/_0041_ ),
    .A2(\adder/norm/_0049_ ),
    .ZN(\adder/norm/_0050_ ));
 NOR2_X1 \adder/norm/_2428_  (.A1(\adder/norm/_0156_ ),
    .A2(\adder/norm/_0090_ ),
    .ZN(\adder/norm/_0052_ ));
 AOI21_X1 \adder/norm/_2429_  (.A(\adder/norm/_0052_ ),
    .B1(\adder/norm/_0048_ ),
    .B2(\adder/norm/_0044_ ),
    .ZN(\adder/norm/_0053_ ));
 NAND2_X1 \adder/norm/_2430_  (.A1(\adder/norm/_0050_ ),
    .A2(\adder/norm/_0053_ ),
    .ZN(\adder/norm/_0054_ ));
 INV_X1 \adder/norm/_2431_  (.A(\adder/norm/_0398_ ),
    .ZN(\adder/norm/_0055_ ));
 XNOR2_X2 \adder/norm/_2432_  (.A(\adder/norm/_0055_ ),
    .B(\adder/norm/_0145_ ),
    .ZN(\adder/norm/_0056_ ));
 XNOR2_X1 \adder/norm/_2433_  (.A(\adder/norm/_0054_ ),
    .B(\adder/norm/_0056_ ),
    .ZN(net68));
 NOR2_X1 \adder/norm/_2434_  (.A1(\adder/norm/_0055_ ),
    .A2(\adder/norm/_0145_ ),
    .ZN(\adder/norm/_0057_ ));
 INV_X1 \adder/norm/_2435_  (.A(\adder/norm/_0056_ ),
    .ZN(\adder/norm/_0058_ ));
 AOI21_X1 \adder/norm/_2436_  (.A(\adder/norm/_0057_ ),
    .B1(\adder/norm/_0054_ ),
    .B2(\adder/norm/_0058_ ),
    .ZN(\adder/norm/_0059_ ));
 INV_X1 \adder/norm/_2437_  (.A(\adder/norm/_0420_ ),
    .ZN(\adder/norm/_0060_ ));
 XNOR2_X1 \adder/norm/_2438_  (.A(\adder/norm/_0060_ ),
    .B(\adder/norm/_0387_ ),
    .ZN(\adder/norm/_0062_ ));
 INV_X1 \adder/norm/_2439_  (.A(\adder/norm/_0062_ ),
    .ZN(\adder/norm/_0063_ ));
 XNOR2_X1 \adder/norm/_2440_  (.A(\adder/norm/_0059_ ),
    .B(\adder/norm/_0063_ ),
    .ZN(net69));
 NOR2_X1 \adder/norm/_2441_  (.A1(\adder/norm/_0056_ ),
    .A2(\adder/norm/_0062_ ),
    .ZN(\adder/norm/_0064_ ));
 NAND2_X1 \adder/norm/_2442_  (.A1(\adder/norm/_0054_ ),
    .A2(\adder/norm/_0064_ ),
    .ZN(\adder/norm/_0065_ ));
 NOR2_X1 \adder/norm/_2443_  (.A1(\adder/norm/_0060_ ),
    .A2(\adder/norm/_0387_ ),
    .ZN(\adder/norm/_0066_ ));
 AOI21_X1 \adder/norm/_2444_  (.A(\adder/norm/_0066_ ),
    .B1(\adder/norm/_0063_ ),
    .B2(\adder/norm/_0057_ ),
    .ZN(\adder/norm/_0067_ ));
 NAND2_X1 \adder/norm/_2445_  (.A1(\adder/norm/_0065_ ),
    .A2(\adder/norm/_0067_ ),
    .ZN(\adder/norm/_0068_ ));
 OAI21_X1 \adder/norm/_2446_  (.A(\adder/norm/_0321_ ),
    .B1(\adder/norm/_0497_ ),
    .B2(\adder/norm/Mant_leadingOne_D[5] ),
    .ZN(\adder/norm/_0069_ ));
 NAND3_X1 \adder/norm/_2447_  (.A1(\adder/norm/_0277_ ),
    .A2(\adder/norm/_0299_ ),
    .A3(\adder/exp_prenorm_d[5] ),
    .ZN(\adder/norm/_0070_ ));
 NAND2_X1 \adder/norm/_2448_  (.A1(\adder/norm/_0069_ ),
    .A2(\adder/norm/_0070_ ),
    .ZN(\adder/norm/_0072_ ));
 XNOR2_X1 \adder/norm/_2449_  (.A(\adder/norm/_0068_ ),
    .B(\adder/norm/_0072_ ),
    .ZN(net70));
 INV_X1 \adder/norm/_2450_  (.A(\adder/norm/_0072_ ),
    .ZN(\adder/norm/_0073_ ));
 NAND2_X1 \adder/norm/_2451_  (.A1(\adder/norm/_0068_ ),
    .A2(\adder/norm/_0073_ ),
    .ZN(\adder/norm/_0074_ ));
 NAND2_X1 \adder/norm/_2452_  (.A1(\adder/norm/_0074_ ),
    .A2(\adder/norm/_0070_ ),
    .ZN(\adder/norm/_0075_ ));
 OAI21_X1 \adder/norm/_2453_  (.A(\adder/norm/_0464_ ),
    .B1(\adder/norm/_0255_ ),
    .B2(\adder/exp_prenorm_d[6] ),
    .ZN(\adder/norm/_0076_ ));
 INV_X1 \adder/norm/_2454_  (.A(\adder/norm/_0076_ ),
    .ZN(\adder/norm/_0077_ ));
 NAND2_X1 \adder/norm/_2455_  (.A1(\adder/norm/_0075_ ),
    .A2(\adder/norm/_0077_ ),
    .ZN(\adder/norm/_0078_ ));
 NAND3_X1 \adder/norm/_2456_  (.A1(\adder/norm/_0074_ ),
    .A2(\adder/norm/_0070_ ),
    .A3(\adder/norm/_0076_ ),
    .ZN(\adder/norm/_0079_ ));
 NAND2_X1 \adder/norm/_2457_  (.A1(\adder/norm/_0078_ ),
    .A2(\adder/norm/_0079_ ),
    .ZN(net72));
 NAND2_X1 \adder/norm/_2458_  (.A1(\adder/norm/_1430_ ),
    .A2(\adder/norm/_0030_ ),
    .ZN(\adder/norm/_0081_ ));
 XNOR2_X1 \adder/norm/_2459_  (.A(\adder/norm/_0081_ ),
    .B(\adder/norm/_1433_ ),
    .ZN(net64));
 NOR2_X4 \adder/norm/_2460_  (.A1(net256),
    .A2(\adder/norm/_0877_ ),
    .ZN(\adder/norm/_0082_ ));
 NAND2_X1 \adder/norm/_2461_  (.A1(net260),
    .A2(\adder/mant_prenorm_d[25] ),
    .ZN(\adder/norm/_0083_ ));
 NAND2_X1 \adder/norm/_2462_  (.A1(\adder/norm/_0083_ ),
    .A2(\adder/norm/_0673_ ),
    .ZN(\adder/norm/_0084_ ));
 TAPCELL_X1 PHY_52 ();
 NAND2_X1 \adder/norm/_2464_  (.A1(net261),
    .A2(\adder/mant_prenorm_d[26] ),
    .ZN(\adder/norm/_0086_ ));
 INV_X1 \adder/norm/_2465_  (.A(\adder/norm/_0086_ ),
    .ZN(\adder/norm/_0087_ ));
 OAI21_X1 \adder/norm/_2466_  (.A(\adder/norm/_0084_ ),
    .B1(\adder/norm/_0673_ ),
    .B2(\adder/norm/_0087_ ),
    .ZN(\adder/norm/_0088_ ));
 OR2_X1 \adder/norm/_2467_  (.A1(\adder/norm/_0088_ ),
    .A2(\adder/norm/_0681_ ),
    .ZN(\adder/norm/_0089_ ));
 TAPCELL_X1 PHY_51 ();
 NAND2_X1 \adder/norm/_2469_  (.A1(net261),
    .A2(\adder/mant_prenorm_d[23] ),
    .ZN(\adder/norm/_0092_ ));
 TAPCELL_X1 PHY_50 ();
 NAND2_X1 \adder/norm/_2471_  (.A1(\adder/norm/_0092_ ),
    .A2(\adder/norm/_0673_ ),
    .ZN(\adder/norm/_0094_ ));
 TAPCELL_X1 PHY_49 ();
 NAND2_X1 \adder/norm/_2473_  (.A1(net261),
    .A2(\adder/mant_prenorm_d[24] ),
    .ZN(\adder/norm/_0096_ ));
 INV_X1 \adder/norm/_2474_  (.A(\adder/norm/_0096_ ),
    .ZN(\adder/norm/_0097_ ));
 OAI21_X1 \adder/norm/_2475_  (.A(\adder/norm/_0094_ ),
    .B1(\adder/norm/_0673_ ),
    .B2(\adder/norm/_0097_ ),
    .ZN(\adder/norm/_0098_ ));
 TAPCELL_X1 PHY_48 ();
 OAI21_X1 \adder/norm/_2477_  (.A(\adder/norm/_0089_ ),
    .B1(\adder/norm/_0098_ ),
    .B2(net82),
    .ZN(\adder/norm/_0100_ ));
 TAPCELL_X1 PHY_47 ();
 NAND2_X1 \adder/norm/_2479_  (.A1(\adder/norm/_0100_ ),
    .A2(\adder/norm/_0694_ ),
    .ZN(\adder/norm/_0103_ ));
 TAPCELL_X1 PHY_46 ();
 NAND2_X1 \adder/norm/_2481_  (.A1(net260),
    .A2(\adder/mant_prenorm_d[21] ),
    .ZN(\adder/norm/_0105_ ));
 NAND2_X1 \adder/norm/_2482_  (.A1(\adder/norm/_0105_ ),
    .A2(\adder/norm/_0673_ ),
    .ZN(\adder/norm/_0106_ ));
 TAPCELL_X1 PHY_45 ();
 TAPCELL_X1 PHY_44 ();
 NAND2_X1 \adder/norm/_2485_  (.A1(net261),
    .A2(\adder/mant_prenorm_d[22] ),
    .ZN(\adder/norm/_0109_ ));
 INV_X1 \adder/norm/_2486_  (.A(\adder/norm/_0109_ ),
    .ZN(\adder/norm/_0110_ ));
 OAI21_X1 \adder/norm/_2487_  (.A(\adder/norm/_0106_ ),
    .B1(\adder/norm/_0673_ ),
    .B2(\adder/norm/_0110_ ),
    .ZN(\adder/norm/_0111_ ));
 NAND2_X1 \adder/norm/_2488_  (.A1(net260),
    .A2(\adder/mant_prenorm_d[20] ),
    .ZN(\adder/norm/_0113_ ));
 NAND2_X1 \adder/norm/_2489_  (.A1(net248),
    .A2(net165),
    .ZN(\adder/norm/_0114_ ));
 MUX2_X1 \adder/norm/_2490_  (.A(\adder/norm/_0113_ ),
    .B(\adder/norm/_0114_ ),
    .S(\adder/norm/_0673_ ),
    .Z(\adder/norm/_0115_ ));
 MUX2_X1 \adder/norm/_2491_  (.A(\adder/norm/_0111_ ),
    .B(\adder/norm/_0115_ ),
    .S(\adder/norm/_0681_ ),
    .Z(\adder/norm/_0116_ ));
 OAI21_X1 \adder/norm/_2492_  (.A(\adder/norm/_0103_ ),
    .B1(\adder/norm/_0116_ ),
    .B2(\adder/norm/_0694_ ),
    .ZN(\adder/norm/_0117_ ));
 TAPCELL_X1 PHY_43 ();
 MUX2_X1 \adder/norm/_2494_  (.A(\adder/norm/_0113_ ),
    .B(\adder/norm/_0105_ ),
    .S(net84),
    .Z(\adder/norm/_0119_ ));
 TAPCELL_X1 PHY_42 ();
 NAND2_X1 \adder/norm/_2496_  (.A1(\adder/norm/_0119_ ),
    .A2(\adder/norm/_0681_ ),
    .ZN(\adder/norm/_0121_ ));
 TAPCELL_X1 PHY_41 ();
 NAND2_X1 \adder/norm/_2498_  (.A1(\adder/norm/_0092_ ),
    .A2(net84),
    .ZN(\adder/norm/_0124_ ));
 TAPCELL_X1 PHY_40 ();
 OAI21_X1 \adder/norm/_2500_  (.A(\adder/norm/_0124_ ),
    .B1(net271),
    .B2(\adder/norm/_0110_ ),
    .ZN(\adder/norm/_0126_ ));
 NAND2_X1 \adder/norm/_2501_  (.A1(\adder/norm/_0126_ ),
    .A2(net82),
    .ZN(\adder/norm/_0127_ ));
 NAND2_X1 \adder/norm/_2502_  (.A1(\adder/norm/_0121_ ),
    .A2(\adder/norm/_0127_ ),
    .ZN(\adder/norm/_0128_ ));
 TAPCELL_X1 PHY_39 ();
 NAND2_X1 \adder/norm/_2504_  (.A1(\adder/norm/_0128_ ),
    .A2(net240),
    .ZN(\adder/norm/_0130_ ));
 NAND2_X1 \adder/norm/_2505_  (.A1(\adder/norm/_0097_ ),
    .A2(\adder/norm/_0673_ ),
    .ZN(\adder/norm/_0131_ ));
 OAI21_X1 \adder/norm/_2506_  (.A(\adder/norm/_0131_ ),
    .B1(\adder/norm/_0673_ ),
    .B2(\adder/norm/_0083_ ),
    .ZN(\adder/norm/_0132_ ));
 NAND2_X1 \adder/norm/_2507_  (.A1(\adder/norm/_0132_ ),
    .A2(\adder/norm/_0681_ ),
    .ZN(\adder/norm/_0133_ ));
 TAPCELL_X1 PHY_38 ();
 NAND2_X1 \adder/norm/_2509_  (.A1(net260),
    .A2(\adder/mant_prenorm_d[27] ),
    .ZN(\adder/norm/_0136_ ));
 NAND2_X1 \adder/norm/_2510_  (.A1(\adder/norm/_0136_ ),
    .A2(net271),
    .ZN(\adder/norm/_0137_ ));
 OAI21_X1 \adder/norm/_2511_  (.A(\adder/norm/_0137_ ),
    .B1(net271),
    .B2(\adder/norm/_0087_ ),
    .ZN(\adder/norm/_0138_ ));
 OAI21_X1 \adder/norm/_2512_  (.A(\adder/norm/_0133_ ),
    .B1(\adder/norm/_0681_ ),
    .B2(\adder/norm/_0138_ ),
    .ZN(\adder/norm/_0139_ ));
 TAPCELL_X1 PHY_37 ();
 OAI21_X1 \adder/norm/_2514_  (.A(\adder/norm/_0130_ ),
    .B1(\adder/norm/_0139_ ),
    .B2(net240),
    .ZN(\adder/norm/_0141_ ));
 INV_X1 \adder/norm/_2515_  (.A(\adder/norm/_0141_ ),
    .ZN(\adder/norm/_0142_ ));
 TAPCELL_X1 PHY_36 ();
 NOR3_X1 \adder/norm/_2517_  (.A1(\adder/norm/_0117_ ),
    .A2(\adder/norm/_0142_ ),
    .A3(net250),
    .ZN(\adder/norm/_0144_ ));
 MUX2_X1 \adder/norm/_2518_  (.A(\adder/norm/_0098_ ),
    .B(\adder/norm/_0111_ ),
    .S(\adder/norm/_0681_ ),
    .Z(\adder/norm/_0146_ ));
 TAPCELL_X1 PHY_35 ();
 TAPCELL_X1 PHY_34 ();
 NAND2_X1 \adder/norm/_2521_  (.A1(\adder/norm/_0126_ ),
    .A2(\adder/norm/_0681_ ),
    .ZN(\adder/norm/_0149_ ));
 TAPCELL_X1 PHY_33 ();
 OAI21_X1 \adder/norm/_2523_  (.A(\adder/norm/_0149_ ),
    .B1(\adder/norm/_0681_ ),
    .B2(\adder/norm/_0132_ ),
    .ZN(\adder/norm/_0151_ ));
 NAND3_X1 \adder/norm/_2524_  (.A1(\adder/norm/_0146_ ),
    .A2(\adder/norm/_0694_ ),
    .A3(\adder/norm/_0151_ ),
    .ZN(\adder/norm/_0152_ ));
 TAPCELL_X1 PHY_32 ();
 NAND2_X1 \adder/norm/_2526_  (.A1(\adder/norm/_0119_ ),
    .A2(net82),
    .ZN(\adder/norm/_0154_ ));
 TAPCELL_X1 PHY_31 ();
 NAND2_X4 \adder/norm/_2528_  (.A1(\adder/norm/_0660_ ),
    .A2(\adder/norm/_1013_ ),
    .ZN(\adder/norm/_0157_ ));
 NOR2_X1 \adder/norm/_2529_  (.A1(\adder/norm/_0157_ ),
    .A2(\adder/norm/_1098_ ),
    .ZN(\adder/norm/_0158_ ));
 NAND2_X1 \adder/norm/_2530_  (.A1(\adder/norm/_0158_ ),
    .A2(\adder/norm/_0673_ ),
    .ZN(\adder/norm/_0159_ ));
 OAI21_X1 \adder/norm/_2531_  (.A(\adder/norm/_0159_ ),
    .B1(\adder/norm/_0673_ ),
    .B2(\adder/norm/_0114_ ),
    .ZN(\adder/norm/_0160_ ));
 OAI21_X1 \adder/norm/_2532_  (.A(\adder/norm/_0154_ ),
    .B1(net82),
    .B2(\adder/norm/_0160_ ),
    .ZN(\adder/norm/_0161_ ));
 NAND2_X1 \adder/norm/_2533_  (.A1(\adder/norm/_0115_ ),
    .A2(net82),
    .ZN(\adder/norm/_0162_ ));
 TAPCELL_X1 PHY_30 ();
 NAND2_X1 \adder/norm/_2535_  (.A1(\adder/norm/_0158_ ),
    .A2(net271),
    .ZN(\adder/norm/_0164_ ));
 NAND2_X1 \adder/norm/_2536_  (.A1(net248),
    .A2(net166),
    .ZN(\adder/norm/_0165_ ));
 OAI21_X1 \adder/norm/_2537_  (.A(\adder/norm/_0164_ ),
    .B1(net271),
    .B2(\adder/norm/_0165_ ),
    .ZN(\adder/norm/_0166_ ));
 OAI21_X1 \adder/norm/_2538_  (.A(\adder/norm/_0162_ ),
    .B1(net82),
    .B2(\adder/norm/_0166_ ),
    .ZN(\adder/norm/_0168_ ));
 NAND2_X1 \adder/norm/_2539_  (.A1(\adder/norm/_0161_ ),
    .A2(\adder/norm/_0168_ ),
    .ZN(\adder/norm/_0169_ ));
 OAI21_X1 \adder/norm/_2540_  (.A(\adder/norm/_0152_ ),
    .B1(\adder/norm/_0694_ ),
    .B2(\adder/norm/_0169_ ),
    .ZN(\adder/norm/_0170_ ));
 NAND3_X1 \adder/norm/_2541_  (.A1(\adder/norm/_0146_ ),
    .A2(net240),
    .A3(\adder/norm/_0151_ ),
    .ZN(\adder/norm/_0171_ ));
 NAND2_X1 \adder/norm/_2542_  (.A1(\adder/norm/_0138_ ),
    .A2(\adder/norm/_0681_ ),
    .ZN(\adder/norm/_0172_ ));
 INV_X1 \adder/norm/_2543_  (.A(\adder/mant_prenorm_d[28] ),
    .ZN(\adder/norm/_0173_ ));
 OAI21_X1 \adder/norm/_2544_  (.A(\adder/norm/_0673_ ),
    .B1(\adder/norm/_0157_ ),
    .B2(\adder/norm/_0173_ ),
    .ZN(\adder/norm/_0174_ ));
 NAND2_X1 \adder/norm/_2545_  (.A1(net261),
    .A2(\adder/mant_prenorm_d[29] ),
    .ZN(\adder/norm/_0175_ ));
 NAND2_X1 \adder/norm/_2546_  (.A1(\adder/norm/_0175_ ),
    .A2(net84),
    .ZN(\adder/norm/_0176_ ));
 NAND2_X1 \adder/norm/_2547_  (.A1(\adder/norm/_0174_ ),
    .A2(\adder/norm/_0176_ ),
    .ZN(\adder/norm/_0177_ ));
 INV_X1 \adder/norm/_2548_  (.A(\adder/norm/_0177_ ),
    .ZN(\adder/norm/_0179_ ));
 OAI21_X1 \adder/norm/_2549_  (.A(\adder/norm/_0172_ ),
    .B1(\adder/norm/_0681_ ),
    .B2(\adder/norm/_0179_ ),
    .ZN(\adder/norm/_0180_ ));
 NAND2_X1 \adder/norm/_2550_  (.A1(\adder/norm/_0088_ ),
    .A2(\adder/norm/_0681_ ),
    .ZN(\adder/norm/_0181_ ));
 NAND3_X1 \adder/norm/_2551_  (.A1(net260),
    .A2(\adder/mant_prenorm_d[28] ),
    .A3(net271),
    .ZN(\adder/norm/_0182_ ));
 OAI21_X1 \adder/norm/_2552_  (.A(\adder/norm/_0182_ ),
    .B1(net271),
    .B2(\adder/norm/_0136_ ),
    .ZN(\adder/norm/_0183_ ));
 OAI21_X1 \adder/norm/_2553_  (.A(\adder/norm/_0181_ ),
    .B1(\adder/norm/_0681_ ),
    .B2(\adder/norm/_0183_ ),
    .ZN(\adder/norm/_0184_ ));
 NAND3_X1 \adder/norm/_2554_  (.A1(\adder/norm/_0180_ ),
    .A2(\adder/norm/_0184_ ),
    .A3(\adder/norm/_0694_ ),
    .ZN(\adder/norm/_0185_ ));
 NAND2_X1 \adder/norm/_2555_  (.A1(\adder/norm/_0171_ ),
    .A2(\adder/norm/_0185_ ),
    .ZN(\adder/norm/_0186_ ));
 NAND3_X1 \adder/norm/_2556_  (.A1(\adder/norm/_0144_ ),
    .A2(\adder/norm/_0170_ ),
    .A3(\adder/norm/_0186_ ),
    .ZN(\adder/norm/_0187_ ));
 AND2_X1 \adder/norm/_2557_  (.A1(net261),
    .A2(\adder/mant_prenorm_d[36] ),
    .ZN(\adder/norm/_0188_ ));
 NAND2_X1 \adder/norm/_2558_  (.A1(\adder/norm/_0188_ ),
    .A2(net271),
    .ZN(\adder/norm/_0190_ ));
 TAPCELL_X1 PHY_29 ();
 NAND2_X1 \adder/norm/_2560_  (.A1(net260),
    .A2(\adder/mant_prenorm_d[35] ),
    .ZN(\adder/norm/_0192_ ));
 OAI21_X1 \adder/norm/_2561_  (.A(\adder/norm/_0190_ ),
    .B1(net271),
    .B2(\adder/norm/_0192_ ),
    .ZN(\adder/norm/_0193_ ));
 TAPCELL_X1 PHY_28 ();
 NAND2_X1 \adder/norm/_2563_  (.A1(\adder/norm/_0193_ ),
    .A2(net82),
    .ZN(\adder/norm/_0195_ ));
 TAPCELL_X1 PHY_27 ();
 NAND2_X1 \adder/norm/_2565_  (.A1(net260),
    .A2(\adder/mant_prenorm_d[33] ),
    .ZN(\adder/norm/_0197_ ));
 NAND2_X1 \adder/norm/_2566_  (.A1(net260),
    .A2(\adder/mant_prenorm_d[34] ),
    .ZN(\adder/norm/_0198_ ));
 MUX2_X1 \adder/norm/_2567_  (.A(\adder/norm/_0197_ ),
    .B(\adder/norm/_0198_ ),
    .S(net271),
    .Z(\adder/norm/_0199_ ));
 OAI21_X1 \adder/norm/_2568_  (.A(\adder/norm/_0195_ ),
    .B1(net82),
    .B2(\adder/norm/_0199_ ),
    .ZN(\adder/norm/_0201_ ));
 NAND2_X1 \adder/norm/_2569_  (.A1(\adder/norm/_0201_ ),
    .A2(\adder/norm/_0694_ ),
    .ZN(\adder/norm/_0202_ ));
 NAND2_X1 \adder/norm/_2570_  (.A1(\adder/norm/_0175_ ),
    .A2(\adder/norm/_0673_ ),
    .ZN(\adder/norm/_0203_ ));
 NAND2_X1 \adder/norm/_2571_  (.A1(net261),
    .A2(\adder/mant_prenorm_d[30] ),
    .ZN(\adder/norm/_0204_ ));
 NAND2_X1 \adder/norm/_2572_  (.A1(\adder/norm/_0204_ ),
    .A2(net84),
    .ZN(\adder/norm/_0205_ ));
 NAND2_X1 \adder/norm/_2573_  (.A1(\adder/norm/_0203_ ),
    .A2(\adder/norm/_0205_ ),
    .ZN(\adder/norm/_0206_ ));
 NAND2_X1 \adder/norm/_2574_  (.A1(\adder/norm/_0206_ ),
    .A2(\adder/norm/_0681_ ),
    .ZN(\adder/norm/_0207_ ));
 NAND3_X1 \adder/norm/_2575_  (.A1(net248),
    .A2(\adder/mant_prenorm_d[32] ),
    .A3(net271),
    .ZN(\adder/norm/_0208_ ));
 NAND2_X1 \adder/norm/_2576_  (.A1(net261),
    .A2(\adder/mant_prenorm_d[31] ),
    .ZN(\adder/norm/_0209_ ));
 OAI21_X1 \adder/norm/_2577_  (.A(\adder/norm/_0208_ ),
    .B1(net271),
    .B2(\adder/norm/_0209_ ),
    .ZN(\adder/norm/_0210_ ));
 OAI21_X1 \adder/norm/_2578_  (.A(\adder/norm/_0207_ ),
    .B1(\adder/norm/_0210_ ),
    .B2(\adder/norm/_0681_ ),
    .ZN(\adder/norm/_0212_ ));
 OAI21_X1 \adder/norm/_2579_  (.A(\adder/norm/_0202_ ),
    .B1(\adder/norm/_0694_ ),
    .B2(\adder/norm/_0212_ ),
    .ZN(\adder/norm/_0213_ ));
 NAND2_X1 \adder/norm/_2580_  (.A1(\adder/norm/_0188_ ),
    .A2(\adder/norm/_0673_ ),
    .ZN(\adder/norm/_0214_ ));
 NAND3_X1 \adder/norm/_2581_  (.A1(net248),
    .A2(\adder/mant_prenorm_d[37] ),
    .A3(net271),
    .ZN(\adder/norm/_0215_ ));
 NAND2_X1 \adder/norm/_2582_  (.A1(\adder/norm/_0214_ ),
    .A2(\adder/norm/_0215_ ),
    .ZN(\adder/norm/_0216_ ));
 NAND2_X1 \adder/norm/_2583_  (.A1(\adder/norm/_0216_ ),
    .A2(net82),
    .ZN(\adder/norm/_0217_ ));
 NAND2_X1 \adder/norm/_2584_  (.A1(\adder/norm/_0198_ ),
    .A2(\adder/norm/_0673_ ),
    .ZN(\adder/norm/_0218_ ));
 NAND2_X1 \adder/norm/_2585_  (.A1(\adder/norm/_0192_ ),
    .A2(net271),
    .ZN(\adder/norm/_0219_ ));
 NAND2_X1 \adder/norm/_2586_  (.A1(\adder/norm/_0218_ ),
    .A2(\adder/norm/_0219_ ),
    .ZN(\adder/norm/_0220_ ));
 OAI21_X1 \adder/norm/_2587_  (.A(\adder/norm/_0217_ ),
    .B1(net82),
    .B2(\adder/norm/_0220_ ),
    .ZN(\adder/norm/_0221_ ));
 NAND3_X1 \adder/norm/_2588_  (.A1(net248),
    .A2(\adder/mant_prenorm_d[33] ),
    .A3(net271),
    .ZN(\adder/norm/_0223_ ));
 NAND2_X1 \adder/norm/_2589_  (.A1(net248),
    .A2(\adder/mant_prenorm_d[32] ),
    .ZN(\adder/norm/_0224_ ));
 OAI21_X1 \adder/norm/_2590_  (.A(\adder/norm/_0223_ ),
    .B1(net84),
    .B2(\adder/norm/_0224_ ),
    .ZN(\adder/norm/_0225_ ));
 NAND2_X1 \adder/norm/_2591_  (.A1(\adder/norm/_0225_ ),
    .A2(net82),
    .ZN(\adder/norm/_0226_ ));
 NAND2_X1 \adder/norm/_2592_  (.A1(\adder/norm/_0204_ ),
    .A2(\adder/norm/_0673_ ),
    .ZN(\adder/norm/_0227_ ));
 NAND2_X1 \adder/norm/_2593_  (.A1(\adder/norm/_0209_ ),
    .A2(net84),
    .ZN(\adder/norm/_0228_ ));
 NAND2_X1 \adder/norm/_2594_  (.A1(\adder/norm/_0227_ ),
    .A2(\adder/norm/_0228_ ),
    .ZN(\adder/norm/_0229_ ));
 OAI21_X1 \adder/norm/_2595_  (.A(\adder/norm/_0226_ ),
    .B1(net82),
    .B2(\adder/norm/_0229_ ),
    .ZN(\adder/norm/_0230_ ));
 MUX2_X1 \adder/norm/_2596_  (.A(\adder/norm/_0221_ ),
    .B(\adder/norm/_0230_ ),
    .S(net240),
    .Z(\adder/norm/_0231_ ));
 OR2_X1 \adder/norm/_2597_  (.A1(\adder/norm/_0212_ ),
    .A2(net240),
    .ZN(\adder/norm/_0232_ ));
 OAI21_X1 \adder/norm/_2598_  (.A(\adder/norm/_0232_ ),
    .B1(\adder/norm/_0694_ ),
    .B2(\adder/norm/_0184_ ),
    .ZN(\adder/norm/_0234_ ));
 NOR3_X1 \adder/norm/_2599_  (.A1(\adder/norm/_0213_ ),
    .A2(\adder/norm/_0231_ ),
    .A3(\adder/norm/_0234_ ),
    .ZN(\adder/norm/_0235_ ));
 NAND2_X1 \adder/norm/_2600_  (.A1(\adder/norm/_0210_ ),
    .A2(\adder/norm/_0681_ ),
    .ZN(\adder/norm/_0236_ ));
 OAI21_X1 \adder/norm/_2601_  (.A(\adder/norm/_0236_ ),
    .B1(\adder/norm/_0199_ ),
    .B2(\adder/norm/_0681_ ),
    .ZN(\adder/norm/_0237_ ));
 NAND2_X1 \adder/norm/_2602_  (.A1(\adder/norm/_0183_ ),
    .A2(\adder/norm/_0681_ ),
    .ZN(\adder/norm/_0238_ ));
 OAI21_X1 \adder/norm/_2603_  (.A(\adder/norm/_0238_ ),
    .B1(\adder/norm/_0681_ ),
    .B2(\adder/norm/_0206_ ),
    .ZN(\adder/norm/_0239_ ));
 MUX2_X1 \adder/norm/_2604_  (.A(\adder/norm/_0237_ ),
    .B(\adder/norm/_0239_ ),
    .S(net240),
    .Z(\adder/norm/_0240_ ));
 NAND2_X1 \adder/norm/_2605_  (.A1(\adder/norm/_0229_ ),
    .A2(net82),
    .ZN(\adder/norm/_0241_ ));
 TAPCELL_X1 PHY_26 ();
 OAI21_X1 \adder/norm/_2607_  (.A(\adder/norm/_0241_ ),
    .B1(net82),
    .B2(\adder/norm/_0179_ ),
    .ZN(\adder/norm/_0243_ ));
 OR2_X1 \adder/norm/_2608_  (.A1(\adder/norm/_0243_ ),
    .A2(\adder/norm/_0694_ ),
    .ZN(\adder/norm/_0245_ ));
 NAND2_X1 \adder/norm/_2609_  (.A1(\adder/norm/_0220_ ),
    .A2(net82),
    .ZN(\adder/norm/_0246_ ));
 OAI21_X1 \adder/norm/_2610_  (.A(\adder/norm/_0246_ ),
    .B1(\adder/norm/_0225_ ),
    .B2(net82),
    .ZN(\adder/norm/_0247_ ));
 OR2_X1 \adder/norm/_2611_  (.A1(\adder/norm/_0247_ ),
    .A2(net240),
    .ZN(\adder/norm/_0248_ ));
 NAND3_X1 \adder/norm/_2612_  (.A1(\adder/norm/_0245_ ),
    .A2(\adder/norm/_0248_ ),
    .A3(net250),
    .ZN(\adder/norm/_0249_ ));
 NAND2_X1 \adder/norm/_2613_  (.A1(\adder/norm/_0230_ ),
    .A2(\adder/norm/_0694_ ),
    .ZN(\adder/norm/_0250_ ));
 OAI21_X1 \adder/norm/_2614_  (.A(\adder/norm/_0250_ ),
    .B1(\adder/norm/_0694_ ),
    .B2(\adder/norm/_0180_ ),
    .ZN(\adder/norm/_0251_ ));
 NOR3_X1 \adder/norm/_2615_  (.A1(\adder/norm/_0240_ ),
    .A2(\adder/norm/_0249_ ),
    .A3(\adder/norm/_0251_ ),
    .ZN(\adder/norm/_0252_ ));
 NAND2_X1 \adder/norm/_2616_  (.A1(\adder/norm/_0235_ ),
    .A2(\adder/norm/_0252_ ),
    .ZN(\adder/norm/_0253_ ));
 NAND2_X1 \adder/norm/_2617_  (.A1(\adder/norm/_0187_ ),
    .A2(\adder/norm/_0253_ ),
    .ZN(\adder/norm/_0254_ ));
 NAND2_X1 \adder/norm/_2618_  (.A1(\adder/norm/_0243_ ),
    .A2(\adder/norm/_0694_ ),
    .ZN(\adder/norm/_0256_ ));
 OAI21_X1 \adder/norm/_2619_  (.A(\adder/norm/_0256_ ),
    .B1(\adder/norm/_0139_ ),
    .B2(\adder/norm/_0694_ ),
    .ZN(\adder/norm/_0257_ ));
 NAND2_X1 \adder/norm/_2620_  (.A1(\adder/norm/_0100_ ),
    .A2(net240),
    .ZN(\adder/norm/_0258_ ));
 NAND2_X1 \adder/norm/_2621_  (.A1(\adder/norm/_0239_ ),
    .A2(\adder/norm/_0694_ ),
    .ZN(\adder/norm/_0259_ ));
 NAND3_X1 \adder/norm/_2622_  (.A1(\adder/norm/_0257_ ),
    .A2(\adder/norm/_0258_ ),
    .A3(\adder/norm/_0259_ ),
    .ZN(\adder/norm/_0260_ ));
 OAI21_X1 \adder/norm/_2623_  (.A(net250),
    .B1(\adder/norm/_0260_ ),
    .B2(\adder/norm/_0117_ ),
    .ZN(\adder/norm/_0261_ ));
 NOR2_X1 \adder/norm/_2624_  (.A1(\adder/norm/_0157_ ),
    .A2(\adder/norm/_0809_ ),
    .ZN(\adder/norm/_0262_ ));
 NAND2_X1 \adder/norm/_2625_  (.A1(\adder/norm/_0262_ ),
    .A2(net271),
    .ZN(\adder/norm/_0263_ ));
 NAND2_X1 \adder/norm/_2626_  (.A1(net248),
    .A2(net167),
    .ZN(\adder/norm/_0264_ ));
 OAI21_X1 \adder/norm/_2627_  (.A(\adder/norm/_0263_ ),
    .B1(net271),
    .B2(\adder/norm/_0264_ ),
    .ZN(\adder/norm/_0265_ ));
 OR2_X1 \adder/norm/_2628_  (.A1(\adder/norm/_0265_ ),
    .A2(net82),
    .ZN(\adder/norm/_0267_ ));
 OAI21_X1 \adder/norm/_2629_  (.A(\adder/norm/_0267_ ),
    .B1(\adder/norm/_0681_ ),
    .B2(\adder/norm/_0166_ ),
    .ZN(\adder/norm/_0268_ ));
 NAND2_X1 \adder/norm/_2630_  (.A1(net248),
    .A2(net168),
    .ZN(\adder/norm/_0269_ ));
 NAND2_X1 \adder/norm/_2631_  (.A1(\adder/norm/_0269_ ),
    .A2(\adder/norm/_0673_ ),
    .ZN(\adder/norm/_0270_ ));
 NOR2_X1 \adder/norm/_2632_  (.A1(\adder/norm/_0157_ ),
    .A2(\adder/norm/_0797_ ),
    .ZN(\adder/norm/_0271_ ));
 OAI21_X1 \adder/norm/_2633_  (.A(\adder/norm/_0270_ ),
    .B1(\adder/norm/_0271_ ),
    .B2(\adder/norm/_0673_ ),
    .ZN(\adder/norm/_0272_ ));
 NAND2_X1 \adder/norm/_2634_  (.A1(\adder/norm/_0272_ ),
    .A2(\adder/norm/_0681_ ),
    .ZN(\adder/norm/_0273_ ));
 NAND2_X1 \adder/norm/_2635_  (.A1(net248),
    .A2(net169),
    .ZN(\adder/norm/_0274_ ));
 NAND2_X1 \adder/norm/_2636_  (.A1(\adder/norm/_0274_ ),
    .A2(\adder/norm/_0673_ ),
    .ZN(\adder/norm/_0275_ ));
 AND2_X1 \adder/norm/_2637_  (.A1(net248),
    .A2(net170),
    .ZN(\adder/norm/_0276_ ));
 OAI21_X1 \adder/norm/_2638_  (.A(\adder/norm/_0275_ ),
    .B1(\adder/norm/_0276_ ),
    .B2(\adder/norm/_0673_ ),
    .ZN(\adder/norm/_0278_ ));
 NAND2_X1 \adder/norm/_2639_  (.A1(\adder/norm/_0278_ ),
    .A2(net82),
    .ZN(\adder/norm/_0279_ ));
 NAND2_X1 \adder/norm/_2640_  (.A1(\adder/norm/_0273_ ),
    .A2(\adder/norm/_0279_ ),
    .ZN(\adder/norm/_0280_ ));
 INV_X1 \adder/norm/_2641_  (.A(\adder/norm/_0280_ ),
    .ZN(\adder/norm/_0281_ ));
 NAND2_X1 \adder/norm/_2642_  (.A1(\adder/norm/_0281_ ),
    .A2(net240),
    .ZN(\adder/norm/_0282_ ));
 NAND2_X1 \adder/norm/_2643_  (.A1(\adder/norm/_0268_ ),
    .A2(\adder/norm/_0282_ ),
    .ZN(\adder/norm/_0283_ ));
 INV_X1 \adder/norm/_2644_  (.A(\adder/norm/_0283_ ),
    .ZN(\adder/norm/_0284_ ));
 OAI21_X1 \adder/norm/_2645_  (.A(\adder/norm/_0284_ ),
    .B1(net240),
    .B2(\adder/norm/_0116_ ),
    .ZN(\adder/norm/_0285_ ));
 NAND3_X1 \adder/norm/_2646_  (.A1(\adder/norm/_0121_ ),
    .A2(\adder/norm/_0694_ ),
    .A3(\adder/norm/_0127_ ),
    .ZN(\adder/norm/_0286_ ));
 NAND2_X1 \adder/norm/_2647_  (.A1(\adder/norm/_0262_ ),
    .A2(\adder/norm/_0673_ ),
    .ZN(\adder/norm/_0287_ ));
 OAI21_X1 \adder/norm/_2648_  (.A(\adder/norm/_0287_ ),
    .B1(\adder/norm/_0673_ ),
    .B2(\adder/norm/_0165_ ),
    .ZN(\adder/norm/_0289_ ));
 OR2_X1 \adder/norm/_2649_  (.A1(\adder/norm/_0289_ ),
    .A2(net82),
    .ZN(\adder/norm/_0290_ ));
 OAI21_X1 \adder/norm/_2650_  (.A(\adder/norm/_0290_ ),
    .B1(\adder/norm/_0681_ ),
    .B2(\adder/norm/_0160_ ),
    .ZN(\adder/norm/_0291_ ));
 OAI21_X1 \adder/norm/_2651_  (.A(\adder/norm/_0286_ ),
    .B1(\adder/norm/_0291_ ),
    .B2(\adder/norm/_0694_ ),
    .ZN(\adder/norm/_0292_ ));
 OAI21_X1 \adder/norm/_2652_  (.A(\adder/norm/_0747_ ),
    .B1(\adder/norm/_0285_ ),
    .B2(\adder/norm/_0292_ ),
    .ZN(\adder/norm/_0293_ ));
 NAND2_X1 \adder/norm/_2653_  (.A1(\adder/norm/_0261_ ),
    .A2(\adder/norm/_0293_ ),
    .ZN(\adder/norm/_0294_ ));
 INV_X1 \adder/norm/_2654_  (.A(\adder/norm/_0294_ ),
    .ZN(\adder/norm/_0295_ ));
 NAND2_X1 \adder/norm/_2655_  (.A1(\adder/norm/_0254_ ),
    .A2(\adder/norm/_0295_ ),
    .ZN(\adder/norm/_0296_ ));
 NAND2_X1 \adder/norm/_2656_  (.A1(net260),
    .A2(\adder/mant_prenorm_d[43] ),
    .ZN(\adder/norm/_0297_ ));
 NAND2_X1 \adder/norm/_2657_  (.A1(\adder/norm/_0297_ ),
    .A2(\adder/norm/_0673_ ),
    .ZN(\adder/norm/_0298_ ));
 AND2_X1 \adder/norm/_2658_  (.A1(net260),
    .A2(\adder/mant_prenorm_d[44] ),
    .ZN(\adder/norm/_0300_ ));
 OAI21_X1 \adder/norm/_2659_  (.A(\adder/norm/_0298_ ),
    .B1(\adder/norm/_0300_ ),
    .B2(\adder/norm/_0673_ ),
    .ZN(\adder/norm/_0301_ ));
 NAND2_X1 \adder/norm/_2660_  (.A1(net260),
    .A2(\adder/mant_prenorm_d[41] ),
    .ZN(\adder/norm/_0302_ ));
 NAND2_X1 \adder/norm/_2661_  (.A1(\adder/norm/_0302_ ),
    .A2(\adder/norm/_0673_ ),
    .ZN(\adder/norm/_0303_ ));
 AND2_X1 \adder/norm/_2662_  (.A1(net261),
    .A2(\adder/mant_prenorm_d[42] ),
    .ZN(\adder/norm/_0304_ ));
 OAI21_X1 \adder/norm/_2663_  (.A(\adder/norm/_0303_ ),
    .B1(\adder/norm/_0304_ ),
    .B2(\adder/norm/_0673_ ),
    .ZN(\adder/norm/_0305_ ));
 MUX2_X1 \adder/norm/_2664_  (.A(\adder/norm/_0301_ ),
    .B(\adder/norm/_0305_ ),
    .S(\adder/norm/_0681_ ),
    .Z(\adder/norm/_0306_ ));
 INV_X1 \adder/norm/_2665_  (.A(\adder/norm/_0306_ ),
    .ZN(\adder/norm/_0307_ ));
 NAND3_X1 \adder/norm/_2666_  (.A1(net248),
    .A2(\adder/mant_prenorm_d[37] ),
    .A3(\adder/norm/_0673_ ),
    .ZN(\adder/norm/_0308_ ));
 NAND2_X1 \adder/norm/_2667_  (.A1(net261),
    .A2(\adder/mant_prenorm_d[38] ),
    .ZN(\adder/norm/_0309_ ));
 OAI21_X1 \adder/norm/_2668_  (.A(\adder/norm/_0308_ ),
    .B1(\adder/norm/_0673_ ),
    .B2(\adder/norm/_0309_ ),
    .ZN(\adder/norm/_0311_ ));
 NAND2_X1 \adder/norm/_2669_  (.A1(\adder/norm/_0311_ ),
    .A2(\adder/norm/_0681_ ),
    .ZN(\adder/norm/_0312_ ));
 NAND2_X1 \adder/norm/_2670_  (.A1(net261),
    .A2(\adder/mant_prenorm_d[39] ),
    .ZN(\adder/norm/_0313_ ));
 NAND2_X1 \adder/norm/_2671_  (.A1(\adder/norm/_0313_ ),
    .A2(\adder/norm/_0673_ ),
    .ZN(\adder/norm/_0314_ ));
 NOR2_X1 \adder/norm/_2672_  (.A1(\adder/norm/_0157_ ),
    .A2(\adder/norm/_0824_ ),
    .ZN(\adder/norm/_0315_ ));
 OAI21_X1 \adder/norm/_2673_  (.A(\adder/norm/_0314_ ),
    .B1(\adder/norm/_0315_ ),
    .B2(\adder/norm/_0673_ ),
    .ZN(\adder/norm/_0316_ ));
 OAI21_X1 \adder/norm/_2674_  (.A(\adder/norm/_0312_ ),
    .B1(\adder/norm/_0681_ ),
    .B2(\adder/norm/_0316_ ),
    .ZN(\adder/norm/_0317_ ));
 OAI22_X1 \adder/norm/_2675_  (.A1(\adder/norm/_0307_ ),
    .A2(\adder/norm/_0716_ ),
    .B1(\adder/norm/_0715_ ),
    .B2(\adder/norm/_0317_ ),
    .ZN(\adder/norm/_0318_ ));
 INV_X1 \adder/norm/_2676_  (.A(\adder/norm/_0318_ ),
    .ZN(\adder/norm/_0319_ ));
 OAI21_X1 \adder/norm/_2677_  (.A(\adder/norm/_0319_ ),
    .B1(net250),
    .B2(\adder/norm/_0213_ ),
    .ZN(\adder/norm/_0320_ ));
 NAND2_X1 \adder/norm/_2678_  (.A1(\adder/norm/_0193_ ),
    .A2(\adder/norm/_0681_ ),
    .ZN(\adder/norm/_0322_ ));
 NAND2_X1 \adder/norm/_2679_  (.A1(\adder/norm/_0311_ ),
    .A2(net82),
    .ZN(\adder/norm/_0323_ ));
 NAND2_X1 \adder/norm/_2680_  (.A1(\adder/norm/_0322_ ),
    .A2(\adder/norm/_0323_ ),
    .ZN(\adder/norm/_0324_ ));
 MUX2_X1 \adder/norm/_2681_  (.A(\adder/norm/_0324_ ),
    .B(\adder/norm/_0237_ ),
    .S(net240),
    .Z(\adder/norm/_0325_ ));
 NAND2_X1 \adder/norm/_2682_  (.A1(\adder/norm/_0309_ ),
    .A2(\adder/norm/_0673_ ),
    .ZN(\adder/norm/_0326_ ));
 NAND2_X1 \adder/norm/_2683_  (.A1(\adder/norm/_0313_ ),
    .A2(net84),
    .ZN(\adder/norm/_0327_ ));
 AND2_X1 \adder/norm/_2684_  (.A1(\adder/norm/_0326_ ),
    .A2(\adder/norm/_0327_ ),
    .ZN(\adder/norm/_0328_ ));
 MUX2_X1 \adder/norm/_2685_  (.A(\adder/norm/_0216_ ),
    .B(\adder/norm/_0328_ ),
    .S(net82),
    .Z(\adder/norm/_0329_ ));
 NAND2_X1 \adder/norm/_2686_  (.A1(\adder/norm/_0329_ ),
    .A2(\adder/norm/_0694_ ),
    .ZN(\adder/norm/_0330_ ));
 OAI21_X1 \adder/norm/_2687_  (.A(\adder/norm/_0330_ ),
    .B1(\adder/norm/_0694_ ),
    .B2(\adder/norm/_0247_ ),
    .ZN(\adder/norm/_0331_ ));
 OAI21_X1 \adder/norm/_2688_  (.A(net250),
    .B1(\adder/norm/_0325_ ),
    .B2(\adder/norm/_0331_ ),
    .ZN(\adder/norm/_0333_ ));
 NAND2_X1 \adder/norm/_2689_  (.A1(\adder/norm/_0320_ ),
    .A2(\adder/norm/_0333_ ),
    .ZN(\adder/norm/_0334_ ));
 NAND2_X1 \adder/norm/_2690_  (.A1(\adder/norm/_0297_ ),
    .A2(net271),
    .ZN(\adder/norm/_0335_ ));
 OAI21_X1 \adder/norm/_2691_  (.A(\adder/norm/_0335_ ),
    .B1(\adder/norm/_0304_ ),
    .B2(net271),
    .ZN(\adder/norm/_0336_ ));
 NAND2_X1 \adder/norm/_2692_  (.A1(net260),
    .A2(\adder/mant_prenorm_d[45] ),
    .ZN(\adder/norm/_0337_ ));
 NAND2_X1 \adder/norm/_2693_  (.A1(\adder/norm/_0337_ ),
    .A2(net271),
    .ZN(\adder/norm/_0338_ ));
 OAI21_X1 \adder/norm/_2694_  (.A(\adder/norm/_0338_ ),
    .B1(\adder/norm/_0300_ ),
    .B2(net271),
    .ZN(\adder/norm/_0339_ ));
 MUX2_X1 \adder/norm/_2695_  (.A(\adder/norm/_0336_ ),
    .B(\adder/norm/_0339_ ),
    .S(net82),
    .Z(\adder/norm/_0340_ ));
 INV_X1 \adder/norm/_2696_  (.A(\adder/norm/_0340_ ),
    .ZN(\adder/norm/_0341_ ));
 NAND2_X1 \adder/norm/_2697_  (.A1(\adder/norm/_0328_ ),
    .A2(\adder/norm/_0681_ ),
    .ZN(\adder/norm/_0342_ ));
 NAND2_X1 \adder/norm/_2698_  (.A1(\adder/norm/_0302_ ),
    .A2(net271),
    .ZN(\adder/norm/_0344_ ));
 OAI21_X1 \adder/norm/_2699_  (.A(\adder/norm/_0344_ ),
    .B1(\adder/norm/_0315_ ),
    .B2(net271),
    .ZN(\adder/norm/_0345_ ));
 OAI21_X1 \adder/norm/_2700_  (.A(\adder/norm/_0342_ ),
    .B1(\adder/norm/_0681_ ),
    .B2(\adder/norm/_0345_ ),
    .ZN(\adder/norm/_0346_ ));
 OAI22_X1 \adder/norm/_2701_  (.A1(\adder/norm/_0341_ ),
    .A2(\adder/norm/_0716_ ),
    .B1(\adder/norm/_0715_ ),
    .B2(\adder/norm/_0346_ ),
    .ZN(\adder/norm/_0347_ ));
 INV_X1 \adder/norm/_2702_  (.A(\adder/norm/_0347_ ),
    .ZN(\adder/norm/_0348_ ));
 TAPCELL_X1 PHY_25 ();
 OAI21_X1 \adder/norm/_2704_  (.A(\adder/norm/_0348_ ),
    .B1(net250),
    .B2(\adder/norm/_0231_ ),
    .ZN(\adder/norm/_0350_ ));
 INV_X1 \adder/norm/_2705_  (.A(\adder/norm/_0350_ ),
    .ZN(\adder/norm/_0351_ ));
 NOR2_X1 \adder/norm/_2706_  (.A1(\adder/norm/_0334_ ),
    .A2(\adder/norm/_0351_ ),
    .ZN(\adder/norm/_0352_ ));
 NAND2_X1 \adder/norm/_2707_  (.A1(\adder/norm/_0260_ ),
    .A2(\adder/norm/_0747_ ),
    .ZN(\adder/norm/_0353_ ));
 NOR2_X1 \adder/norm/_2708_  (.A1(\adder/norm/_0251_ ),
    .A2(net250),
    .ZN(\adder/norm/_0355_ ));
 OAI22_X1 \adder/norm/_2709_  (.A1(\adder/norm/_0716_ ),
    .A2(\adder/norm/_0346_ ),
    .B1(\adder/norm/_0221_ ),
    .B2(\adder/norm/_0715_ ),
    .ZN(\adder/norm/_0356_ ));
 OAI21_X1 \adder/norm/_2710_  (.A(\adder/norm/_0353_ ),
    .B1(\adder/norm/_0355_ ),
    .B2(\adder/norm/_0356_ ),
    .ZN(\adder/norm/_0357_ ));
 OR2_X1 \adder/norm/_2711_  (.A1(\adder/norm/_0305_ ),
    .A2(\adder/norm/_0681_ ),
    .ZN(\adder/norm/_0358_ ));
 OAI21_X1 \adder/norm/_2712_  (.A(\adder/norm/_0358_ ),
    .B1(net82),
    .B2(\adder/norm/_0316_ ),
    .ZN(\adder/norm/_0359_ ));
 OAI22_X1 \adder/norm/_2713_  (.A1(\adder/norm/_0359_ ),
    .A2(\adder/norm/_0716_ ),
    .B1(\adder/norm/_0324_ ),
    .B2(\adder/norm/_0715_ ),
    .ZN(\adder/norm/_0360_ ));
 INV_X1 \adder/norm/_2714_  (.A(\adder/norm/_0360_ ),
    .ZN(\adder/norm/_0361_ ));
 OAI21_X1 \adder/norm/_2715_  (.A(\adder/norm/_0361_ ),
    .B1(\adder/norm/_0240_ ),
    .B2(net250),
    .ZN(\adder/norm/_0362_ ));
 OAI22_X1 \adder/norm/_2716_  (.A1(\adder/norm/_0201_ ),
    .A2(\adder/norm/_0715_ ),
    .B1(\adder/norm/_0317_ ),
    .B2(\adder/norm/_0716_ ),
    .ZN(\adder/norm/_0363_ ));
 INV_X1 \adder/norm/_2717_  (.A(\adder/norm/_0363_ ),
    .ZN(\adder/norm/_0364_ ));
 OAI21_X1 \adder/norm/_2718_  (.A(\adder/norm/_0364_ ),
    .B1(\adder/norm/_0234_ ),
    .B2(net250),
    .ZN(\adder/norm/_0366_ ));
 NAND2_X1 \adder/norm/_2719_  (.A1(\adder/norm/_0362_ ),
    .A2(\adder/norm/_0366_ ),
    .ZN(\adder/norm/_0367_ ));
 NOR2_X1 \adder/norm/_2720_  (.A1(\adder/norm/_0357_ ),
    .A2(\adder/norm/_0367_ ),
    .ZN(\adder/norm/_0368_ ));
 NAND2_X1 \adder/norm/_2721_  (.A1(\adder/norm/_0352_ ),
    .A2(\adder/norm/_0368_ ),
    .ZN(\adder/norm/_0369_ ));
 NOR2_X1 \adder/norm/_2722_  (.A1(\adder/norm/_0296_ ),
    .A2(\adder/norm/_0369_ ),
    .ZN(\adder/norm/_0370_ ));
 NOR2_X1 \adder/norm/_2723_  (.A1(\adder/norm/_0325_ ),
    .A2(net250),
    .ZN(\adder/norm/_0371_ ));
 NAND2_X1 \adder/norm/_2724_  (.A1(net248),
    .A2(\adder/mant_prenorm_d[46] ),
    .ZN(\adder/norm/_0372_ ));
 MUX2_X1 \adder/norm/_2725_  (.A(\adder/norm/_0372_ ),
    .B(\adder/norm/_0337_ ),
    .S(\adder/norm/_0673_ ),
    .Z(\adder/norm/_0373_ ));
 MUX2_X1 \adder/norm/_2726_  (.A(\adder/norm/_0301_ ),
    .B(\adder/norm/_0373_ ),
    .S(net82),
    .Z(\adder/norm/_0374_ ));
 INV_X1 \adder/norm/_2727_  (.A(\adder/norm/_0374_ ),
    .ZN(\adder/norm/_0375_ ));
 OAI22_X1 \adder/norm/_2728_  (.A1(\adder/norm/_0375_ ),
    .A2(\adder/norm/_0716_ ),
    .B1(\adder/norm/_0359_ ),
    .B2(\adder/norm/_0715_ ),
    .ZN(\adder/norm/_0377_ ));
 NOR2_X1 \adder/norm/_2729_  (.A1(\adder/norm/_0331_ ),
    .A2(net250),
    .ZN(\adder/norm/_0378_ ));
 OR2_X1 \adder/norm/_2730_  (.A1(\adder/norm/_0336_ ),
    .A2(\adder/norm/_0681_ ),
    .ZN(\adder/norm/_0379_ ));
 OAI21_X1 \adder/norm/_2731_  (.A(\adder/norm/_0379_ ),
    .B1(net82),
    .B2(\adder/norm/_0345_ ),
    .ZN(\adder/norm/_0380_ ));
 NAND2_X1 \adder/norm/_2732_  (.A1(\adder/norm/_0339_ ),
    .A2(\adder/norm/_0681_ ),
    .ZN(\adder/norm/_0381_ ));
 OAI22_X1 \adder/norm/_2733_  (.A1(\adder/norm/_0372_ ),
    .A2(net271),
    .B1(\adder/norm/_0861_ ),
    .B2(\adder/norm/_0877_ ),
    .ZN(\adder/norm/_0382_ ));
 OAI21_X1 \adder/norm/_2734_  (.A(\adder/norm/_0381_ ),
    .B1(\adder/norm/_0681_ ),
    .B2(\adder/norm/_0382_ ),
    .ZN(\adder/norm/_0383_ ));
 INV_X1 \adder/norm/_2735_  (.A(\adder/norm/_0383_ ),
    .ZN(\adder/norm/_0384_ ));
 OAI22_X1 \adder/norm/_2736_  (.A1(\adder/norm/_0380_ ),
    .A2(\adder/norm/_0715_ ),
    .B1(\adder/norm/_0384_ ),
    .B2(\adder/norm/_0716_ ),
    .ZN(\adder/norm/_0385_ ));
 OAI22_X1 \adder/norm/_2737_  (.A1(\adder/norm/_0371_ ),
    .A2(\adder/norm/_0377_ ),
    .B1(\adder/norm/_0378_ ),
    .B2(\adder/norm/_0385_ ),
    .ZN(\adder/norm/_0386_ ));
 NAND2_X1 \adder/norm/_2738_  (.A1(\adder/norm/_0141_ ),
    .A2(net250),
    .ZN(\adder/norm/_0388_ ));
 NAND2_X1 \adder/norm/_2739_  (.A1(\adder/norm/_0264_ ),
    .A2(net84),
    .ZN(\adder/norm/_0389_ ));
 OAI21_X1 \adder/norm/_2740_  (.A(\adder/norm/_0389_ ),
    .B1(\adder/norm/_0276_ ),
    .B2(net271),
    .ZN(\adder/norm/_0390_ ));
 NAND2_X1 \adder/norm/_2741_  (.A1(\adder/norm/_0390_ ),
    .A2(net82),
    .ZN(\adder/norm/_0391_ ));
 NAND2_X1 \adder/norm/_2742_  (.A1(\adder/norm/_0271_ ),
    .A2(\adder/norm/_0673_ ),
    .ZN(\adder/norm/_0392_ ));
 OAI21_X1 \adder/norm/_2743_  (.A(\adder/norm/_0392_ ),
    .B1(\adder/norm/_0673_ ),
    .B2(\adder/norm/_0274_ ),
    .ZN(\adder/norm/_0393_ ));
 OAI21_X1 \adder/norm/_2744_  (.A(\adder/norm/_0391_ ),
    .B1(\adder/norm/_0393_ ),
    .B2(net82),
    .ZN(\adder/norm/_0394_ ));
 OR2_X1 \adder/norm/_2745_  (.A1(\adder/norm/_0394_ ),
    .A2(\adder/norm/_0694_ ),
    .ZN(\adder/norm/_0395_ ));
 OAI21_X1 \adder/norm/_2746_  (.A(\adder/norm/_0395_ ),
    .B1(\adder/norm/_0291_ ),
    .B2(net240),
    .ZN(\adder/norm/_0396_ ));
 OAI21_X1 \adder/norm/_2747_  (.A(\adder/norm/_0388_ ),
    .B1(\adder/norm/_0396_ ),
    .B2(net250),
    .ZN(\adder/norm/_0397_ ));
 AND3_X1 \adder/norm/_2748_  (.A1(\adder/norm/_0245_ ),
    .A2(\adder/norm/_0248_ ),
    .A3(\adder/norm/_0747_ ),
    .ZN(\adder/norm/_0399_ ));
 OAI22_X1 \adder/norm/_2749_  (.A1(\adder/norm/_0380_ ),
    .A2(\adder/norm/_0716_ ),
    .B1(\adder/norm/_0329_ ),
    .B2(\adder/norm/_0715_ ),
    .ZN(\adder/norm/_0400_ ));
 OAI21_X1 \adder/norm/_2750_  (.A(\adder/norm/_0397_ ),
    .B1(\adder/norm/_0399_ ),
    .B2(\adder/norm/_0400_ ),
    .ZN(\adder/norm/_0401_ ));
 NAND2_X1 \adder/norm/_2751_  (.A1(net248),
    .A2(net171),
    .ZN(\adder/norm/_0402_ ));
 NAND2_X1 \adder/norm/_2752_  (.A1(\adder/norm/_0402_ ),
    .A2(\adder/norm/_0673_ ),
    .ZN(\adder/norm/_0403_ ));
 NOR2_X1 \adder/norm/_2753_  (.A1(\adder/norm/_0157_ ),
    .A2(\adder/norm/_0784_ ),
    .ZN(\adder/norm/_0404_ ));
 OAI21_X1 \adder/norm/_2754_  (.A(\adder/norm/_0403_ ),
    .B1(\adder/norm/_0673_ ),
    .B2(\adder/norm/_0404_ ),
    .ZN(\adder/norm/_0405_ ));
 NAND2_X1 \adder/norm/_2755_  (.A1(\adder/norm/_0405_ ),
    .A2(\adder/norm/_0681_ ),
    .ZN(\adder/norm/_0406_ ));
 AND2_X1 \adder/norm/_2756_  (.A1(net248),
    .A2(net172),
    .ZN(\adder/norm/_0407_ ));
 NAND2_X1 \adder/norm/_2757_  (.A1(\adder/norm/_0407_ ),
    .A2(net83),
    .ZN(\adder/norm/_0408_ ));
 NAND2_X1 \adder/norm/_2758_  (.A1(net248),
    .A2(net173),
    .ZN(\adder/norm/_0410_ ));
 OAI21_X1 \adder/norm/_2759_  (.A(\adder/norm/_0408_ ),
    .B1(net83),
    .B2(\adder/norm/_0410_ ),
    .ZN(\adder/norm/_0411_ ));
 OAI21_X1 \adder/norm/_2760_  (.A(\adder/norm/_0406_ ),
    .B1(\adder/norm/_0411_ ),
    .B2(\adder/norm/_0681_ ),
    .ZN(\adder/norm/_0412_ ));
 NAND2_X1 \adder/norm/_2761_  (.A1(\adder/norm/_0412_ ),
    .A2(net240),
    .ZN(\adder/norm/_0413_ ));
 OAI21_X1 \adder/norm/_2762_  (.A(\adder/norm/_0413_ ),
    .B1(net240),
    .B2(\adder/norm/_0281_ ),
    .ZN(\adder/norm/_0414_ ));
 OAI21_X1 \adder/norm/_2763_  (.A(\adder/norm/_0673_ ),
    .B1(\adder/norm/_0157_ ),
    .B2(\adder/norm/_0770_ ),
    .ZN(\adder/norm/_0415_ ));
 AND2_X1 \adder/norm/_2764_  (.A1(net248),
    .A2(net174),
    .ZN(\adder/norm/_0416_ ));
 OAI21_X1 \adder/norm/_2765_  (.A(\adder/norm/_0415_ ),
    .B1(\adder/norm/_0416_ ),
    .B2(\adder/norm/_0673_ ),
    .ZN(\adder/norm/_0417_ ));
 NAND2_X1 \adder/norm/_2766_  (.A1(\adder/norm/_0417_ ),
    .A2(\adder/norm/_0681_ ),
    .ZN(\adder/norm/_0418_ ));
 NAND3_X1 \adder/norm/_2767_  (.A1(net248),
    .A2(net175),
    .A3(net83),
    .ZN(\adder/norm/_0419_ ));
 NAND2_X1 \adder/norm/_2768_  (.A1(net248),
    .A2(net176),
    .ZN(\adder/norm/_0421_ ));
 OAI21_X1 \adder/norm/_2769_  (.A(\adder/norm/_0419_ ),
    .B1(net83),
    .B2(\adder/norm/_0421_ ),
    .ZN(\adder/norm/_0422_ ));
 OAI21_X1 \adder/norm/_2770_  (.A(\adder/norm/_0418_ ),
    .B1(\adder/norm/_0681_ ),
    .B2(\adder/norm/_0422_ ),
    .ZN(\adder/norm/_0423_ ));
 NAND2_X1 \adder/norm/_2771_  (.A1(\adder/norm/_0423_ ),
    .A2(\adder/norm/_0694_ ),
    .ZN(\adder/norm/_0424_ ));
 NAND2_X1 \adder/norm/_2772_  (.A1(net248),
    .A2(net177),
    .ZN(\adder/norm/_0425_ ));
 NAND2_X1 \adder/norm/_2773_  (.A1(\adder/norm/_0425_ ),
    .A2(\adder/norm/_0673_ ),
    .ZN(\adder/norm/_0426_ ));
 NAND2_X1 \adder/norm/_2774_  (.A1(net248),
    .A2(net178),
    .ZN(\adder/norm/_0427_ ));
 NAND2_X1 \adder/norm/_2775_  (.A1(\adder/norm/_0427_ ),
    .A2(net83),
    .ZN(\adder/norm/_0428_ ));
 NAND3_X1 \adder/norm/_2776_  (.A1(\adder/norm/_0426_ ),
    .A2(\adder/norm/_0428_ ),
    .A3(net81),
    .ZN(\adder/norm/_0429_ ));
 NOR3_X1 \adder/norm/_2777_  (.A1(\adder/norm/_0157_ ),
    .A2(\adder/norm/_0878_ ),
    .A3(\adder/norm/_0673_ ),
    .ZN(\adder/norm/_0430_ ));
 NAND2_X1 \adder/norm/_2778_  (.A1(\adder/norm/_0430_ ),
    .A2(\adder/norm/_0681_ ),
    .ZN(\adder/norm/_0432_ ));
 NAND2_X1 \adder/norm/_2779_  (.A1(\adder/norm/_0429_ ),
    .A2(\adder/norm/_0432_ ),
    .ZN(\adder/norm/_0433_ ));
 OAI21_X1 \adder/norm/_2780_  (.A(\adder/norm/_0424_ ),
    .B1(\adder/norm/_0694_ ),
    .B2(\adder/norm/_0433_ ),
    .ZN(\adder/norm/_0434_ ));
 MUX2_X1 \adder/norm/_2781_  (.A(\adder/norm/_0414_ ),
    .B(\adder/norm/_0434_ ),
    .S(\adder/norm/_0747_ ),
    .Z(\adder/norm/_0435_ ));
 NAND3_X1 \adder/norm/_2782_  (.A1(net248),
    .A2(net179),
    .A3(\adder/norm/_0673_ ),
    .ZN(\adder/norm/_0436_ ));
 OAI21_X1 \adder/norm/_2783_  (.A(\adder/norm/_0436_ ),
    .B1(\adder/norm/_0673_ ),
    .B2(\adder/norm/_0402_ ),
    .ZN(\adder/norm/_0437_ ));
 NAND2_X1 \adder/norm/_2784_  (.A1(\adder/norm/_0437_ ),
    .A2(net81),
    .ZN(\adder/norm/_0438_ ));
 NAND2_X1 \adder/norm/_2785_  (.A1(\adder/norm/_0421_ ),
    .A2(net83),
    .ZN(\adder/norm/_0439_ ));
 OAI21_X1 \adder/norm/_2786_  (.A(\adder/norm/_0439_ ),
    .B1(\adder/norm/_0416_ ),
    .B2(net83),
    .ZN(\adder/norm/_0440_ ));
 OAI21_X1 \adder/norm/_2787_  (.A(\adder/norm/_0438_ ),
    .B1(net81),
    .B2(\adder/norm/_0440_ ),
    .ZN(\adder/norm/_0441_ ));
 OR2_X1 \adder/norm/_2788_  (.A1(\adder/norm/_0441_ ),
    .A2(\adder/norm/_0694_ ),
    .ZN(\adder/norm/_0443_ ));
 NAND2_X1 \adder/norm/_2789_  (.A1(\adder/norm/_0410_ ),
    .A2(net83),
    .ZN(\adder/norm/_0444_ ));
 OAI21_X1 \adder/norm/_2790_  (.A(\adder/norm/_0444_ ),
    .B1(net83),
    .B2(\adder/norm/_0404_ ),
    .ZN(\adder/norm/_0445_ ));
 INV_X1 \adder/norm/_2791_  (.A(\adder/norm/_0445_ ),
    .ZN(\adder/norm/_0446_ ));
 NAND2_X1 \adder/norm/_2792_  (.A1(\adder/norm/_0446_ ),
    .A2(\adder/norm/_0681_ ),
    .ZN(\adder/norm/_0447_ ));
 NAND2_X1 \adder/norm/_2793_  (.A1(\adder/norm/_0269_ ),
    .A2(net83),
    .ZN(\adder/norm/_0448_ ));
 OAI21_X1 \adder/norm/_2794_  (.A(\adder/norm/_0448_ ),
    .B1(\adder/norm/_0407_ ),
    .B2(net83),
    .ZN(\adder/norm/_0449_ ));
 OAI21_X1 \adder/norm/_2795_  (.A(\adder/norm/_0447_ ),
    .B1(\adder/norm/_0681_ ),
    .B2(\adder/norm/_0449_ ),
    .ZN(\adder/norm/_0450_ ));
 OAI21_X1 \adder/norm/_2796_  (.A(\adder/norm/_0443_ ),
    .B1(net240),
    .B2(\adder/norm/_0450_ ),
    .ZN(\adder/norm/_0451_ ));
 NAND2_X1 \adder/norm/_2797_  (.A1(\adder/norm/_0451_ ),
    .A2(net250),
    .ZN(\adder/norm/_0452_ ));
 NAND3_X1 \adder/norm/_2798_  (.A1(net248),
    .A2(net180),
    .A3(\adder/norm/_0673_ ),
    .ZN(\adder/norm/_0454_ ));
 OAI21_X1 \adder/norm/_2799_  (.A(\adder/norm/_0454_ ),
    .B1(\adder/norm/_0673_ ),
    .B2(\adder/norm/_0425_ ),
    .ZN(\adder/norm/_0455_ ));
 NAND2_X1 \adder/norm/_2800_  (.A1(\adder/norm/_0455_ ),
    .A2(\adder/norm/_0681_ ),
    .ZN(\adder/norm/_0456_ ));
 NAND3_X1 \adder/norm/_2801_  (.A1(net248),
    .A2(net181),
    .A3(net83),
    .ZN(\adder/norm/_0457_ ));
 OAI21_X1 \adder/norm/_2802_  (.A(\adder/norm/_0457_ ),
    .B1(net83),
    .B2(\adder/norm/_0427_ ),
    .ZN(\adder/norm/_0458_ ));
 INV_X1 \adder/norm/_2803_  (.A(\adder/norm/_0458_ ),
    .ZN(\adder/norm/_0459_ ));
 OAI21_X1 \adder/norm/_2804_  (.A(\adder/norm/_0456_ ),
    .B1(\adder/norm/_0681_ ),
    .B2(\adder/norm/_0459_ ),
    .ZN(\adder/norm/_0460_ ));
 NAND2_X1 \adder/norm/_2805_  (.A1(\adder/norm/_0460_ ),
    .A2(\adder/norm/_0694_ ),
    .ZN(\adder/norm/_0461_ ));
 INV_X1 \adder/norm/_2806_  (.A(\adder/norm/_0461_ ),
    .ZN(\adder/norm/_0462_ ));
 OAI21_X1 \adder/norm/_2807_  (.A(\adder/norm/_0452_ ),
    .B1(net250),
    .B2(\adder/norm/_0462_ ),
    .ZN(\adder/norm/_0463_ ));
 NAND2_X1 \adder/norm/_2808_  (.A1(\adder/norm/_0435_ ),
    .A2(\adder/norm/_0463_ ),
    .ZN(\adder/norm/_0465_ ));
 NOR3_X1 \adder/norm/_2809_  (.A1(\adder/norm/_0386_ ),
    .A2(\adder/norm/_0401_ ),
    .A3(\adder/norm/_0465_ ),
    .ZN(\adder/norm/_0466_ ));
 NAND2_X1 \adder/norm/_2810_  (.A1(\adder/norm/_0370_ ),
    .A2(\adder/norm/_0466_ ),
    .ZN(\adder/norm/_0467_ ));
 NAND2_X1 \adder/norm/_2811_  (.A1(\adder/norm/_0289_ ),
    .A2(net82),
    .ZN(\adder/norm/_0468_ ));
 OAI21_X1 \adder/norm/_2812_  (.A(\adder/norm/_0468_ ),
    .B1(net82),
    .B2(\adder/norm/_0390_ ),
    .ZN(\adder/norm/_0469_ ));
 NAND2_X1 \adder/norm/_2813_  (.A1(\adder/norm/_0265_ ),
    .A2(net82),
    .ZN(\adder/norm/_0470_ ));
 OAI21_X1 \adder/norm/_2814_  (.A(\adder/norm/_0470_ ),
    .B1(net82),
    .B2(\adder/norm/_0278_ ),
    .ZN(\adder/norm/_0471_ ));
 NOR2_X1 \adder/norm/_2815_  (.A1(\adder/norm/_0469_ ),
    .A2(\adder/norm/_0471_ ),
    .ZN(\adder/norm/_0472_ ));
 NAND2_X1 \adder/norm/_2816_  (.A1(\adder/norm/_0472_ ),
    .A2(\adder/norm/_0694_ ),
    .ZN(\adder/norm/_0473_ ));
 NAND2_X1 \adder/norm/_2817_  (.A1(\adder/norm/_0449_ ),
    .A2(\adder/norm/_0681_ ),
    .ZN(\adder/norm/_0474_ ));
 OAI21_X1 \adder/norm/_2818_  (.A(\adder/norm/_0474_ ),
    .B1(\adder/norm/_0393_ ),
    .B2(\adder/norm/_0681_ ),
    .ZN(\adder/norm/_0476_ ));
 NAND2_X1 \adder/norm/_2819_  (.A1(\adder/norm/_0272_ ),
    .A2(net82),
    .ZN(\adder/norm/_0477_ ));
 OAI21_X1 \adder/norm/_2820_  (.A(\adder/norm/_0477_ ),
    .B1(\adder/norm/_0411_ ),
    .B2(net82),
    .ZN(\adder/norm/_0478_ ));
 NAND2_X1 \adder/norm/_2821_  (.A1(\adder/norm/_0476_ ),
    .A2(\adder/norm/_0478_ ),
    .ZN(\adder/norm/_0479_ ));
 OAI21_X1 \adder/norm/_2822_  (.A(\adder/norm/_0473_ ),
    .B1(\adder/norm/_0694_ ),
    .B2(\adder/norm/_0479_ ),
    .ZN(\adder/norm/_0480_ ));
 NAND2_X1 \adder/norm/_2823_  (.A1(\adder/norm/_0472_ ),
    .A2(net240),
    .ZN(\adder/norm/_0481_ ));
 OAI21_X1 \adder/norm/_2824_  (.A(\adder/norm/_0481_ ),
    .B1(net240),
    .B2(\adder/norm/_0169_ ),
    .ZN(\adder/norm/_0482_ ));
 NAND2_X1 \adder/norm/_2825_  (.A1(\adder/norm/_0480_ ),
    .A2(\adder/norm/_0482_ ),
    .ZN(\adder/norm/_0483_ ));
 NOR2_X1 \adder/norm/_2826_  (.A1(\adder/norm/_0483_ ),
    .A2(\adder/norm/_0285_ ),
    .ZN(\adder/norm/_0484_ ));
 NOR3_X1 \adder/norm/_2827_  (.A1(\adder/norm/_0396_ ),
    .A2(\adder/norm/_0292_ ),
    .A3(\adder/norm/_0747_ ),
    .ZN(\adder/norm/_0485_ ));
 NAND2_X1 \adder/norm/_2828_  (.A1(\adder/norm/_0484_ ),
    .A2(\adder/norm/_0485_ ),
    .ZN(\adder/norm/_0487_ ));
 NAND2_X1 \adder/norm/_2829_  (.A1(\adder/norm/_0445_ ),
    .A2(net81),
    .ZN(\adder/norm/_0488_ ));
 OAI21_X1 \adder/norm/_2830_  (.A(\adder/norm/_0488_ ),
    .B1(\adder/norm/_0437_ ),
    .B2(net81),
    .ZN(\adder/norm/_0489_ ));
 NAND2_X1 \adder/norm/_2831_  (.A1(\adder/norm/_0405_ ),
    .A2(net81),
    .ZN(\adder/norm/_0490_ ));
 OAI21_X1 \adder/norm/_2832_  (.A(\adder/norm/_0490_ ),
    .B1(net81),
    .B2(\adder/norm/_0422_ ),
    .ZN(\adder/norm/_0491_ ));
 NAND2_X1 \adder/norm/_2833_  (.A1(\adder/norm/_0489_ ),
    .A2(\adder/norm/_0491_ ),
    .ZN(\adder/norm/_0492_ ));
 AND2_X1 \adder/norm/_2834_  (.A1(\adder/norm/_0417_ ),
    .A2(net81),
    .ZN(\adder/norm/_0493_ ));
 AOI21_X1 \adder/norm/_2835_  (.A(net81),
    .B1(\adder/norm/_0426_ ),
    .B2(\adder/norm/_0428_ ),
    .ZN(\adder/norm/_0494_ ));
 AOI22_X1 \adder/norm/_2836_  (.A1(\adder/norm/_0493_ ),
    .A2(\adder/norm/_0440_ ),
    .B1(\adder/norm/_0459_ ),
    .B2(\adder/norm/_0494_ ),
    .ZN(\adder/norm/_0495_ ));
 MUX2_X1 \adder/norm/_2837_  (.A(\adder/norm/_0492_ ),
    .B(\adder/norm/_0495_ ),
    .S(net240),
    .Z(\adder/norm/_0496_ ));
 INV_X1 \adder/norm/_2838_  (.A(\adder/norm/_0496_ ),
    .ZN(\adder/norm/_0498_ ));
 OR2_X1 \adder/norm/_2839_  (.A1(\adder/norm/_0412_ ),
    .A2(net240),
    .ZN(\adder/norm/_0499_ ));
 OAI21_X1 \adder/norm/_2840_  (.A(\adder/norm/_0499_ ),
    .B1(\adder/norm/_0694_ ),
    .B2(\adder/norm/_0423_ ),
    .ZN(\adder/norm/_0500_ ));
 NOR2_X1 \adder/norm/_2841_  (.A1(\adder/norm/_0500_ ),
    .A2(net250),
    .ZN(\adder/norm/_0501_ ));
 AND2_X1 \adder/norm/_2842_  (.A1(\adder/norm/_0451_ ),
    .A2(\adder/norm/_0414_ ),
    .ZN(\adder/norm/_0502_ ));
 NAND3_X1 \adder/norm/_2843_  (.A1(\adder/norm/_0498_ ),
    .A2(\adder/norm/_0501_ ),
    .A3(\adder/norm/_0502_ ),
    .ZN(\adder/norm/_0503_ ));
 NAND2_X1 \adder/norm/_2844_  (.A1(\adder/norm/_0394_ ),
    .A2(\adder/norm/_0694_ ),
    .ZN(\adder/norm/_0504_ ));
 OAI21_X1 \adder/norm/_2845_  (.A(\adder/norm/_0504_ ),
    .B1(\adder/norm/_0694_ ),
    .B2(\adder/norm/_0450_ ),
    .ZN(\adder/norm/_0505_ ));
 NOR2_X1 \adder/norm/_2846_  (.A1(\adder/norm/_0479_ ),
    .A2(net240),
    .ZN(\adder/norm/_0506_ ));
 NOR2_X1 \adder/norm/_2847_  (.A1(\adder/norm/_0492_ ),
    .A2(\adder/norm/_0694_ ),
    .ZN(\adder/norm/_0507_ ));
 OAI21_X1 \adder/norm/_2848_  (.A(\adder/norm/_0505_ ),
    .B1(\adder/norm/_0506_ ),
    .B2(\adder/norm/_0507_ ),
    .ZN(\adder/norm/_0509_ ));
 OAI21_X1 \adder/norm/_2849_  (.A(\adder/norm/_0487_ ),
    .B1(\adder/norm/_0503_ ),
    .B2(\adder/norm/_0509_ ),
    .ZN(\adder/norm/_0510_ ));
 NAND3_X1 \adder/norm/_2850_  (.A1(\adder/norm/_0171_ ),
    .A2(net250),
    .A3(\adder/norm/_0185_ ),
    .ZN(\adder/norm/_0511_ ));
 OAI21_X1 \adder/norm/_2851_  (.A(\adder/norm/_0511_ ),
    .B1(\adder/norm/_0482_ ),
    .B2(net250),
    .ZN(\adder/norm/_0512_ ));
 NOR2_X1 \adder/norm/_2852_  (.A1(\adder/norm/_0480_ ),
    .A2(net250),
    .ZN(\adder/norm/_0513_ ));
 NOR2_X1 \adder/norm/_2853_  (.A1(\adder/norm/_0170_ ),
    .A2(\adder/norm/_0747_ ),
    .ZN(\adder/norm/_0514_ ));
 NOR3_X1 \adder/norm/_2854_  (.A1(\adder/norm/_0512_ ),
    .A2(\adder/norm/_0513_ ),
    .A3(\adder/norm/_0514_ ),
    .ZN(\adder/norm/_0515_ ));
 NAND2_X1 \adder/norm/_2855_  (.A1(\adder/norm/_0510_ ),
    .A2(\adder/norm/_0515_ ),
    .ZN(\adder/norm/_0516_ ));
 OAI21_X1 \adder/norm/_2856_  (.A(\adder/norm/_0889_ ),
    .B1(\adder/norm/_0467_ ),
    .B2(\adder/norm/_0516_ ),
    .ZN(\adder/norm/_0517_ ));
 AND2_X1 \adder/norm/_2857_  (.A1(\adder/norm/_0295_ ),
    .A2(\adder/norm/_0397_ ),
    .ZN(\adder/norm/_0518_ ));
 NAND3_X1 \adder/norm/_2858_  (.A1(\adder/norm/_0510_ ),
    .A2(\adder/norm/_0518_ ),
    .A3(\adder/norm/_0515_ ),
    .ZN(\adder/norm/_0520_ ));
 NAND2_X1 \adder/norm/_2859_  (.A1(\adder/norm/_0520_ ),
    .A2(\adder/norm/_0870_ ),
    .ZN(\adder/norm/_0521_ ));
 AOI22_X1 \adder/norm/_2860_  (.A1(\adder/norm/_0435_ ),
    .A2(\adder/norm/_0463_ ),
    .B1(\adder/norm/_0760_ ),
    .B2(\adder/norm/_0869_ ),
    .ZN(\adder/norm/_0522_ ));
 NAND2_X1 \adder/norm/_2861_  (.A1(\adder/norm/_0441_ ),
    .A2(\adder/norm/_0694_ ),
    .ZN(\adder/norm/_0523_ ));
 NAND2_X1 \adder/norm/_2862_  (.A1(\adder/norm/_0460_ ),
    .A2(net240),
    .ZN(\adder/norm/_0524_ ));
 NAND2_X1 \adder/norm/_2863_  (.A1(\adder/norm/_0433_ ),
    .A2(\adder/norm/_0694_ ),
    .ZN(\adder/norm/_0525_ ));
 NAND3_X1 \adder/norm/_2864_  (.A1(\adder/norm/_0523_ ),
    .A2(\adder/norm/_0524_ ),
    .A3(\adder/norm/_0525_ ),
    .ZN(\adder/norm/_0526_ ));
 OR2_X1 \adder/norm/_2865_  (.A1(\adder/norm/_0455_ ),
    .A2(\adder/norm/_0430_ ),
    .ZN(\adder/norm/_0527_ ));
 NAND3_X1 \adder/norm/_2866_  (.A1(\adder/norm/_0527_ ),
    .A2(\adder/norm/_0694_ ),
    .A3(net81),
    .ZN(\adder/norm/_0528_ ));
 INV_X1 \adder/norm/_2867_  (.A(\adder/norm/_0528_ ),
    .ZN(\adder/norm/_0529_ ));
 AOI21_X1 \adder/norm/_2868_  (.A(\adder/norm/_0526_ ),
    .B1(\adder/norm/_0747_ ),
    .B2(\adder/norm/_0529_ ),
    .ZN(\adder/norm/_0531_ ));
 NAND2_X1 \adder/norm/_2869_  (.A1(\adder/norm/_0495_ ),
    .A2(\adder/norm/_0694_ ),
    .ZN(\adder/norm/_0532_ ));
 NAND2_X1 \adder/norm/_2870_  (.A1(\adder/norm/_0527_ ),
    .A2(net81),
    .ZN(\adder/norm/_0533_ ));
 OAI21_X1 \adder/norm/_2871_  (.A(\adder/norm/_0532_ ),
    .B1(\adder/norm/_0694_ ),
    .B2(\adder/norm/_0533_ ),
    .ZN(\adder/norm/_0534_ ));
 INV_X1 \adder/norm/_2872_  (.A(\adder/norm/_0534_ ),
    .ZN(\adder/norm/_0535_ ));
 OAI21_X1 \adder/norm/_2873_  (.A(\adder/norm/_0531_ ),
    .B1(\adder/norm/_0535_ ),
    .B2(net250),
    .ZN(\adder/norm/_0536_ ));
 NOR2_X1 \adder/norm/_2874_  (.A1(\adder/norm/_0498_ ),
    .A2(\adder/norm/_0747_ ),
    .ZN(\adder/norm/_0537_ ));
 NOR2_X1 \adder/norm/_2875_  (.A1(\adder/norm/_0536_ ),
    .A2(\adder/norm/_0537_ ),
    .ZN(\adder/norm/_0538_ ));
 NOR3_X1 \adder/norm/_2876_  (.A1(\adder/norm/_0500_ ),
    .A2(\adder/norm/_0462_ ),
    .A3(\adder/norm/_0529_ ),
    .ZN(\adder/norm/_0539_ ));
 NAND2_X1 \adder/norm/_2877_  (.A1(\adder/norm/_0539_ ),
    .A2(\adder/norm/_0535_ ),
    .ZN(\adder/norm/_0540_ ));
 NAND2_X1 \adder/norm/_2878_  (.A1(\adder/norm/_0540_ ),
    .A2(net250),
    .ZN(\adder/norm/_0542_ ));
 INV_X1 \adder/norm/_2879_  (.A(\adder/norm/_0509_ ),
    .ZN(\adder/norm/_0543_ ));
 NAND2_X1 \adder/norm/_2880_  (.A1(\adder/norm/_0543_ ),
    .A2(\adder/norm/_0434_ ),
    .ZN(\adder/norm/_0544_ ));
 NAND2_X1 \adder/norm/_2881_  (.A1(\adder/norm/_0544_ ),
    .A2(net250),
    .ZN(\adder/norm/_0545_ ));
 NAND3_X1 \adder/norm/_2882_  (.A1(\adder/norm/_0538_ ),
    .A2(\adder/norm/_0542_ ),
    .A3(\adder/norm/_0545_ ),
    .ZN(\adder/norm/_0546_ ));
 AOI21_X1 \adder/norm/_2883_  (.A(\adder/norm/_0522_ ),
    .B1(\adder/norm/_0546_ ),
    .B2(\adder/norm/_1372_ ),
    .ZN(\adder/norm/_0547_ ));
 NAND2_X1 \adder/norm/_2884_  (.A1(\adder/norm/_0521_ ),
    .A2(\adder/norm/_0547_ ),
    .ZN(\adder/norm/_0548_ ));
 INV_X1 \adder/norm/_2885_  (.A(\adder/norm/_0548_ ),
    .ZN(\adder/norm/_0549_ ));
 NAND2_X1 \adder/norm/_2886_  (.A1(\adder/norm/_0517_ ),
    .A2(\adder/norm/_0549_ ),
    .ZN(\adder/norm/_0550_ ));
 NOR3_X1 \adder/norm/_2887_  (.A1(\adder/norm/_0716_ ),
    .A2(\adder/norm/_0681_ ),
    .A3(\adder/norm/_0673_ ),
    .ZN(\adder/norm/_0551_ ));
 NOR2_X1 \adder/norm/_2888_  (.A1(\adder/norm/_1372_ ),
    .A2(\adder/norm/_0551_ ),
    .ZN(\adder/norm/_0553_ ));
 NOR3_X1 \adder/norm/_2889_  (.A1(\adder/norm/_1068_ ),
    .A2(net256),
    .A3(\adder/norm/_0553_ ),
    .ZN(\adder/norm/_0554_ ));
 NAND2_X1 \adder/norm/_2890_  (.A1(\adder/norm/_0550_ ),
    .A2(\adder/norm/_0554_ ),
    .ZN(\adder/norm/_0555_ ));
 AND3_X1 \adder/norm/_2891_  (.A1(\adder/norm/_1067_ ),
    .A2(\adder/norm/_0889_ ),
    .A3(\adder/norm/_0551_ ),
    .ZN(\adder/norm/_0556_ ));
 AOI22_X1 \adder/norm/_2892_  (.A1(\adder/norm/_0556_ ),
    .A2(\adder/norm/_0660_ ),
    .B1(\adder/norm/_0656_ ),
    .B2(\adder/norm/_0653_ ),
    .ZN(\adder/norm/_0557_ ));
 NAND2_X1 \adder/norm/_2893_  (.A1(\adder/norm/_0555_ ),
    .A2(\adder/norm/_0557_ ),
    .ZN(\adder/norm/_0558_ ));
 NOR4_X1 \adder/norm/_2894_  (.A1(net182),
    .A2(net183),
    .A3(net184),
    .A4(net185),
    .ZN(\adder/norm/_0559_ ));
 NOR4_X1 \adder/norm/_2895_  (.A1(net186),
    .A2(net187),
    .A3(net188),
    .A4(net189),
    .ZN(\adder/norm/_0560_ ));
 NOR4_X1 \adder/norm/_2896_  (.A1(net190),
    .A2(net191),
    .A3(net192),
    .A4(net193),
    .ZN(\adder/norm/_0561_ ));
 NOR4_X1 \adder/norm/_2897_  (.A1(net194),
    .A2(net195),
    .A3(net196),
    .A4(net197),
    .ZN(\adder/norm/_0562_ ));
 NAND4_X1 \adder/norm/_2898_  (.A1(\adder/norm/_0559_ ),
    .A2(\adder/norm/_0560_ ),
    .A3(\adder/norm/_0561_ ),
    .A4(\adder/norm/_0562_ ),
    .ZN(\adder/norm/_0564_ ));
 NOR4_X1 \adder/norm/_2899_  (.A1(net198),
    .A2(net199),
    .A3(net200),
    .A4(net201),
    .ZN(\adder/norm/_0565_ ));
 NOR4_X1 \adder/norm/_2900_  (.A1(\adder/mant_prenorm_d[23] ),
    .A2(\adder/mant_prenorm_d[22] ),
    .A3(\adder/mant_prenorm_d[21] ),
    .A4(\adder/mant_prenorm_d[20] ),
    .ZN(\adder/norm/_0566_ ));
 NOR4_X1 \adder/norm/_2901_  (.A1(\adder/mant_prenorm_d[27] ),
    .A2(\adder/mant_prenorm_d[26] ),
    .A3(\adder/mant_prenorm_d[25] ),
    .A4(\adder/mant_prenorm_d[24] ),
    .ZN(\adder/norm/_0567_ ));
 NOR4_X1 \adder/norm/_2902_  (.A1(\adder/mant_prenorm_d[31] ),
    .A2(\adder/mant_prenorm_d[30] ),
    .A3(\adder/mant_prenorm_d[29] ),
    .A4(\adder/mant_prenorm_d[28] ),
    .ZN(\adder/norm/_0568_ ));
 NAND4_X1 \adder/norm/_2903_  (.A1(\adder/norm/_0565_ ),
    .A2(\adder/norm/_0566_ ),
    .A3(\adder/norm/_0567_ ),
    .A4(\adder/norm/_0568_ ),
    .ZN(\adder/norm/_0569_ ));
 NOR4_X1 \adder/norm/_2904_  (.A1(\adder/mant_prenorm_d[35] ),
    .A2(\adder/mant_prenorm_d[34] ),
    .A3(\adder/mant_prenorm_d[33] ),
    .A4(\adder/mant_prenorm_d[32] ),
    .ZN(\adder/norm/_0570_ ));
 NOR4_X1 \adder/norm/_2905_  (.A1(\adder/mant_prenorm_d[46] ),
    .A2(\adder/mant_prenorm_d[47] ),
    .A3(\adder/mant_prenorm_d[45] ),
    .A4(\adder/mant_prenorm_d[44] ),
    .ZN(\adder/norm/_0571_ ));
 NOR4_X1 \adder/norm/_2906_  (.A1(\adder/mant_prenorm_d[39] ),
    .A2(\adder/mant_prenorm_d[38] ),
    .A3(\adder/mant_prenorm_d[37] ),
    .A4(\adder/mant_prenorm_d[36] ),
    .ZN(\adder/norm/_0572_ ));
 NOR4_X1 \adder/norm/_2907_  (.A1(\adder/mant_prenorm_d[43] ),
    .A2(\adder/mant_prenorm_d[42] ),
    .A3(\adder/mant_prenorm_d[41] ),
    .A4(\adder/mant_prenorm_d[40] ),
    .ZN(\adder/norm/_0573_ ));
 NAND4_X1 \adder/norm/_2908_  (.A1(\adder/norm/_0570_ ),
    .A2(\adder/norm/_0571_ ),
    .A3(\adder/norm/_0572_ ),
    .A4(\adder/norm/_0573_ ),
    .ZN(\adder/norm/_0575_ ));
 OR4_X1 \adder/norm/_2909_  (.A1(\adder/norm/_0557_ ),
    .A2(\adder/norm/_0564_ ),
    .A3(\adder/norm/_0569_ ),
    .A4(\adder/norm/_0575_ ),
    .ZN(\adder/norm/_0576_ ));
 NAND2_X1 \adder/norm/_2910_  (.A1(\adder/norm/_0558_ ),
    .A2(\adder/norm/_0576_ ),
    .ZN(\adder/norm/_0577_ ));
 AOI22_X1 \adder/norm/_2911_  (.A1(\adder/norm/_0851_ ),
    .A2(\adder/norm/_0868_ ),
    .B1(\adder/norm/_1261_ ),
    .B2(\adder/norm/_1264_ ),
    .ZN(\adder/norm/_0578_ ));
 NAND2_X1 \adder/norm/_2912_  (.A1(\adder/norm/_0989_ ),
    .A2(\adder/norm/_1005_ ),
    .ZN(\adder/norm/_0579_ ));
 AND4_X1 \adder/norm/_2913_  (.A1(\adder/norm/_0643_ ),
    .A2(\adder/norm/_0578_ ),
    .A3(\adder/norm/_0757_ ),
    .A4(\adder/norm/_0579_ ),
    .ZN(\adder/norm/_0580_ ));
 AOI22_X1 \adder/norm/_2914_  (.A1(\adder/norm/_0750_ ),
    .A2(\adder/norm/_0720_ ),
    .B1(\adder/norm/_1247_ ),
    .B2(\adder/norm/_1250_ ),
    .ZN(\adder/norm/_0581_ ));
 AOI21_X1 \adder/norm/_2915_  (.A(\adder/norm/_0759_ ),
    .B1(\adder/norm/_0918_ ),
    .B2(\adder/norm/_0936_ ),
    .ZN(\adder/norm/_0582_ ));
 AND2_X1 \adder/norm/_2916_  (.A1(\adder/norm/_0581_ ),
    .A2(\adder/norm/_0582_ ),
    .ZN(\adder/norm/_0583_ ));
 OAI21_X1 \adder/norm/_2917_  (.A(\adder/norm/_0754_ ),
    .B1(\adder/norm/_0580_ ),
    .B2(\adder/norm/_0583_ ),
    .ZN(\adder/norm/_0584_ ));
 NAND2_X1 \adder/norm/_2918_  (.A1(\adder/norm/_0796_ ),
    .A2(\adder/norm/_0819_ ),
    .ZN(\adder/norm/_0586_ ));
 NAND2_X1 \adder/norm/_2919_  (.A1(\adder/norm/_0953_ ),
    .A2(\adder/norm/_0971_ ),
    .ZN(\adder/norm/_0587_ ));
 NAND2_X1 \adder/norm/_2920_  (.A1(\adder/norm/_1254_ ),
    .A2(\adder/norm/_1257_ ),
    .ZN(\adder/norm/_0588_ ));
 NAND4_X1 \adder/norm/_2921_  (.A1(\adder/norm/_0586_ ),
    .A2(\adder/norm/_0587_ ),
    .A3(\adder/norm/_0588_ ),
    .A4(\adder/norm/_0761_ ),
    .ZN(\adder/norm/_0589_ ));
 NAND2_X1 \adder/norm/_2922_  (.A1(\adder/norm/_1010_ ),
    .A2(\adder/norm/_0820_ ),
    .ZN(\adder/norm/_0590_ ));
 OR3_X1 \adder/norm/_2923_  (.A1(\adder/norm/_1268_ ),
    .A2(\adder/norm/_0887_ ),
    .A3(\adder/norm/_0590_ ),
    .ZN(\adder/norm/_0591_ ));
 NAND4_X1 \adder/norm/_2924_  (.A1(\adder/norm/_0584_ ),
    .A2(\adder/norm/_1067_ ),
    .A3(\adder/norm/_0589_ ),
    .A4(\adder/norm/_0591_ ),
    .ZN(\adder/norm/_0592_ ));
 NAND2_X1 \adder/norm/_2925_  (.A1(\adder/norm/_0577_ ),
    .A2(\adder/norm/_0592_ ),
    .ZN(\adder/norm/_0593_ ));
 INV_X1 \adder/norm/_2926_  (.A(\adder/norm/_1310_ ),
    .ZN(\adder/norm/_0594_ ));
 NAND3_X1 \adder/norm/_2927_  (.A1(\adder/norm/_0593_ ),
    .A2(\adder/norm/_1320_ ),
    .A3(\adder/norm/_0594_ ),
    .ZN(\adder/norm/_0595_ ));
 INV_X1 \adder/norm/_2928_  (.A(\adder/norm/_1320_ ),
    .ZN(\adder/norm/_0597_ ));
 NAND2_X1 \adder/norm/_2929_  (.A1(\adder/norm/_0597_ ),
    .A2(\adder/norm/_1310_ ),
    .ZN(\adder/norm/_0598_ ));
 NAND2_X1 \adder/norm/_2930_  (.A1(\adder/norm/_0595_ ),
    .A2(\adder/norm/_0598_ ),
    .ZN(net49));
 NOR2_X1 \adder/norm/_2931_  (.A1(\adder/norm/_0594_ ),
    .A2(\adder/norm/_0597_ ),
    .ZN(\adder/norm/_0599_ ));
 XOR2_X1 \adder/norm/_2932_  (.A(\adder/norm/_0599_ ),
    .B(\adder/norm/_1292_ ),
    .Z(net60));
 XNOR2_X1 \adder/norm/_2933_  (.A(\adder/norm/_1321_ ),
    .B(\adder/norm/_1356_ ),
    .ZN(net71));
 INV_X1 \adder/norm/_2934_  (.A(\adder/norm/_1321_ ),
    .ZN(\adder/norm/_0600_ ));
 AOI21_X1 \adder/norm/_2935_  (.A(\adder/norm/_1339_ ),
    .B1(\adder/norm/_0600_ ),
    .B2(\adder/norm/_1356_ ),
    .ZN(\adder/norm/_0601_ ));
 NOR2_X1 \adder/norm/_2936_  (.A1(\adder/norm/_0601_ ),
    .A2(\adder/norm/_1358_ ),
    .ZN(net74));
 XOR2_X1 \adder/norm/_2937_  (.A(\adder/norm/_1358_ ),
    .B(\adder/norm/_1394_ ),
    .Z(net75));
 NAND2_X1 \adder/norm/_2938_  (.A1(\adder/norm/_1358_ ),
    .A2(\adder/norm/_1394_ ),
    .ZN(\adder/norm/_0603_ ));
 XNOR2_X1 \adder/norm/_2939_  (.A(\adder/norm/_0603_ ),
    .B(\adder/norm/_1377_ ),
    .ZN(net76));
 NAND3_X1 \adder/norm/_2940_  (.A1(\adder/norm/_1358_ ),
    .A2(\adder/norm/_1394_ ),
    .A3(\adder/norm/_1377_ ),
    .ZN(\adder/norm/_0604_ ));
 XNOR2_X1 \adder/norm/_2941_  (.A(\adder/norm/_0604_ ),
    .B(\adder/norm/_1426_ ),
    .ZN(net77));
 NAND4_X2 \adder/norm/_2942_  (.A1(\adder/norm/_1358_ ),
    .A2(\adder/norm/_1426_ ),
    .A3(\adder/norm/_1394_ ),
    .A4(\adder/norm/_1377_ ),
    .ZN(\adder/norm/_0605_ ));
 XNOR2_X1 \adder/norm/_2943_  (.A(\adder/norm/_0605_ ),
    .B(\adder/norm/_1410_ ),
    .ZN(net78));
 XNOR2_X1 \adder/norm/_2944_  (.A(\adder/norm/_1429_ ),
    .B(\adder/norm/_1209_ ),
    .ZN(net79));
 INV_X1 \adder/norm/_2945_  (.A(\adder/norm/_1410_ ),
    .ZN(\adder/norm/_0606_ ));
 NOR2_X1 \adder/norm/_2946_  (.A1(\adder/norm/_0605_ ),
    .A2(\adder/norm/_0606_ ),
    .ZN(\adder/norm/_0607_ ));
 AOI21_X1 \adder/norm/_2947_  (.A(\adder/norm/_1171_ ),
    .B1(\adder/norm/_0607_ ),
    .B2(\adder/norm/_1209_ ),
    .ZN(\adder/norm/_0608_ ));
 INV_X1 \adder/norm/_2948_  (.A(\adder/norm/_1210_ ),
    .ZN(\adder/norm/_0610_ ));
 AOI21_X1 \adder/norm/_2949_  (.A(\adder/norm/_0608_ ),
    .B1(\adder/norm/_0607_ ),
    .B2(\adder/norm/_0610_ ),
    .ZN(net80));
 AND3_X1 \adder/norm/_2950_  (.A1(\adder/norm/_0607_ ),
    .A2(\adder/norm/_0610_ ),
    .A3(\adder/norm/_1074_ ),
    .ZN(\adder/norm/_0611_ ));
 AOI21_X1 \adder/norm/_2951_  (.A(\adder/norm/_1074_ ),
    .B1(\adder/norm/_0607_ ),
    .B2(\adder/norm/_0610_ ),
    .ZN(\adder/norm/_0612_ ));
 NOR2_X1 \adder/norm/_2952_  (.A1(\adder/norm/_0611_ ),
    .A2(\adder/norm/_0612_ ),
    .ZN(net50));
 AOI21_X1 \adder/norm/_2953_  (.A(\adder/norm/_0611_ ),
    .B1(\adder/norm/_1116_ ),
    .B2(\adder/norm/_1132_ ),
    .ZN(\adder/norm/_0613_ ));
 AOI21_X1 \adder/norm/_2954_  (.A(\adder/norm/_0613_ ),
    .B1(\adder/norm/_0607_ ),
    .B2(\adder/norm/_1211_ ),
    .ZN(net51));
 NAND3_X1 \adder/norm/_2955_  (.A1(\adder/norm/_1358_ ),
    .A2(\adder/norm/_1428_ ),
    .A3(\adder/norm/_1211_ ),
    .ZN(\adder/norm/_0614_ ));
 XOR2_X1 \adder/norm/_2956_  (.A(\adder/norm/_0614_ ),
    .B(\adder/norm/_1015_ ),
    .Z(net52));
 NOR2_X1 \adder/norm/_2957_  (.A1(\adder/norm/_0614_ ),
    .A2(\adder/norm/_1015_ ),
    .ZN(\adder/norm/_0615_ ));
 XNOR2_X1 \adder/norm/_2958_  (.A(\adder/norm/_0615_ ),
    .B(\adder/norm/_0896_ ),
    .ZN(net53));
 NOR3_X1 \adder/norm/_2959_  (.A1(\adder/norm/_0614_ ),
    .A2(\adder/norm/_1015_ ),
    .A3(\adder/norm/_0896_ ),
    .ZN(\adder/norm/_0617_ ));
 XNOR2_X1 \adder/norm/_2960_  (.A(\adder/norm/_0617_ ),
    .B(\adder/norm/_1271_ ),
    .ZN(net54));
 NAND3_X1 \adder/norm/_2961_  (.A1(\adder/norm/_0617_ ),
    .A2(\adder/norm/_1266_ ),
    .A3(\adder/norm/_1270_ ),
    .ZN(\adder/norm/_0618_ ));
 XOR2_X1 \adder/norm/_2962_  (.A(\adder/norm/_0618_ ),
    .B(\adder/norm/_1244_ ),
    .Z(net55));
 XNOR2_X1 \adder/norm/_2963_  (.A(\adder/norm/_1430_ ),
    .B(\adder/norm/_0008_ ),
    .ZN(net56));
 INV_X1 \adder/norm/_2964_  (.A(\adder/norm/_1430_ ),
    .ZN(\adder/norm/_0619_ ));
 NOR2_X1 \adder/norm/_2965_  (.A1(\adder/norm/_0619_ ),
    .A2(\adder/norm/_0008_ ),
    .ZN(\adder/norm/_0620_ ));
 XNOR2_X1 \adder/norm/_2966_  (.A(\adder/norm/_0620_ ),
    .B(\adder/norm/_0000_ ),
    .ZN(net57));
 NAND2_X1 \adder/norm/_2967_  (.A1(\adder/norm/_1430_ ),
    .A2(\adder/norm/_0009_ ),
    .ZN(\adder/norm/_0621_ ));
 XOR2_X1 \adder/norm/_2968_  (.A(\adder/norm/_0621_ ),
    .B(\adder/norm/_0027_ ),
    .Z(net58));
 NOR2_X1 \adder/norm/_2969_  (.A1(\adder/norm/_0621_ ),
    .A2(\adder/norm/_0027_ ),
    .ZN(\adder/norm/_0623_ ));
 XNOR2_X1 \adder/norm/_2970_  (.A(\adder/norm/_0623_ ),
    .B(\adder/norm/_0018_ ),
    .ZN(net59));
 NOR2_X1 \adder/norm/_2971_  (.A1(\adder/norm/_0619_ ),
    .A2(\adder/norm/_0029_ ),
    .ZN(\adder/norm/_0624_ ));
 XNOR2_X1 \adder/norm/_2972_  (.A(\adder/norm/_0624_ ),
    .B(\adder/norm/_1465_ ),
    .ZN(net61));
 NOR3_X1 \adder/norm/_2973_  (.A1(\adder/norm/_0619_ ),
    .A2(\adder/norm/_1465_ ),
    .A3(\adder/norm/_0029_ ),
    .ZN(\adder/norm/_0625_ ));
 XNOR2_X1 \adder/norm/_2974_  (.A(\adder/norm/_0625_ ),
    .B(\adder/norm/_1457_ ),
    .ZN(net62));
 NAND2_X1 \adder/norm/_2975_  (.A1(\adder/norm/_0624_ ),
    .A2(\adder/norm/_1466_ ),
    .ZN(\adder/norm/_0626_ ));
 INV_X1 \adder/norm/_2976_  (.A(\adder/norm/_1449_ ),
    .ZN(\adder/norm/_0627_ ));
 XNOR2_X1 \adder/norm/_2977_  (.A(\adder/norm/_0626_ ),
    .B(\adder/norm/_0627_ ),
    .ZN(net63));
 NAND3_X1 \adder/norm/_2978_  (.A1(\adder/norm/_0624_ ),
    .A2(\adder/norm/_0627_ ),
    .A3(\adder/norm/_1466_ ),
    .ZN(\adder/norm/_0629_ ));
 INV_X1 \adder/norm/_2979_  (.A(\adder/norm/_1441_ ),
    .ZN(\adder/norm/_0630_ ));
 OR2_X1 \adder/norm/_2980_  (.A1(\adder/norm/_0629_ ),
    .A2(\adder/norm/_0630_ ),
    .ZN(\adder/norm/_0631_ ));
 NAND2_X1 \adder/norm/_2981_  (.A1(\adder/norm/_0629_ ),
    .A2(\adder/norm/_0630_ ),
    .ZN(\adder/norm/_0632_ ));
 NAND3_X1 \adder/norm/_2982_  (.A1(\adder/norm/_1430_ ),
    .A2(\adder/norm/_0646_ ),
    .A3(\adder/norm/_0030_ ),
    .ZN(\adder/norm/_0633_ ));
 NAND3_X1 \adder/norm/_2983_  (.A1(\adder/norm/_0631_ ),
    .A2(\adder/norm/_0632_ ),
    .A3(\adder/norm/_0633_ ),
    .ZN(\adder/mant_norm_d[23] ));
 INV_X1 \converter/_162_  (.A(net3),
    .ZN(\converter/_095_ ));
 INV_X1 \converter/_163_  (.A(net2),
    .ZN(\converter/_096_ ));
 NAND2_X1 \converter/_164_  (.A1(\converter/_095_ ),
    .A2(\converter/_096_ ),
    .ZN(\converter/_097_ ));
 TAPCELL_X1 PHY_24 ();
 NOR4_X4 \converter/_166_  (.A1(\converter/_097_ ),
    .A2(net5),
    .A3(net4),
    .A4(net6),
    .ZN(\converter/_099_ ));
 INV_X4 \converter/_167_  (.A(\converter/_099_ ),
    .ZN(\converter/_100_ ));
 TAPCELL_X1 PHY_23 ();
 TAPCELL_X1 PHY_22 ();
 NAND2_X1 \converter/_170_  (.A1(\converter/_100_ ),
    .A2(net1),
    .ZN(\converter/_103_ ));
 INV_X1 \converter/_171_  (.A(\converter/_103_ ),
    .ZN(\operand_fp16_fp32[13] ));
 INV_X1 \converter/_172_  (.A(net16),
    .ZN(\converter/_104_ ));
 INV_X2 \converter/_173_  (.A(net14),
    .ZN(\converter/_105_ ));
 TAPCELL_X1 PHY_21 ();
 OAI21_X1 \converter/_175_  (.A(\converter/_104_ ),
    .B1(\converter/_105_ ),
    .B2(net15),
    .ZN(\converter/_107_ ));
 NOR2_X4 \converter/_176_  (.A1(net16),
    .A2(net15),
    .ZN(\converter/_108_ ));
 NOR2_X4 \converter/_177_  (.A1(net14),
    .A2(net13),
    .ZN(\converter/_109_ ));
 NAND2_X4 \converter/_178_  (.A1(\converter/_108_ ),
    .A2(\converter/_109_ ),
    .ZN(\converter/_110_ ));
 INV_X4 \converter/_179_  (.A(\converter/_110_ ),
    .ZN(\converter/_111_ ));
 INV_X2 \converter/_180_  (.A(net12),
    .ZN(\converter/_112_ ));
 TAPCELL_X1 PHY_20 ();
 INV_X1 \converter/_182_  (.A(net10),
    .ZN(\converter/_114_ ));
 TAPCELL_X1 PHY_19 ();
 OAI21_X2 \converter/_184_  (.A(\converter/_112_ ),
    .B1(\converter/_114_ ),
    .B2(net11),
    .ZN(\converter/_116_ ));
 AOI21_X4 \converter/_185_  (.A(\converter/_107_ ),
    .B1(\converter/_111_ ),
    .B2(\converter/_116_ ),
    .ZN(\converter/_117_ ));
 NOR2_X1 \converter/_186_  (.A1(net12),
    .A2(net11),
    .ZN(\converter/_118_ ));
 NOR2_X1 \converter/_187_  (.A1(net10),
    .A2(net9),
    .ZN(\converter/_119_ ));
 NAND2_X2 \converter/_188_  (.A1(\converter/_118_ ),
    .A2(\converter/_119_ ),
    .ZN(\converter/_120_ ));
 NOR2_X4 \converter/_189_  (.A1(\converter/_120_ ),
    .A2(\converter/_110_ ),
    .ZN(\converter/_121_ ));
 INV_X1 \converter/_190_  (.A(net8),
    .ZN(\converter/_122_ ));
 NAND2_X1 \converter/_191_  (.A1(\converter/_122_ ),
    .A2(net1),
    .ZN(\converter/_123_ ));
 NAND2_X4 \converter/_192_  (.A1(\converter/_121_ ),
    .A2(\converter/_123_ ),
    .ZN(\converter/_124_ ));
 NAND2_X4 \converter/_193_  (.A1(\converter/_124_ ),
    .A2(\converter/_117_ ),
    .ZN(\converter/_125_ ));
 INV_X4 \converter/_194_  (.A(net262),
    .ZN(\converter/_126_ ));
 INV_X2 \converter/_195_  (.A(\converter/_120_ ),
    .ZN(\converter/_127_ ));
 NAND2_X1 \converter/_196_  (.A1(\converter/_127_ ),
    .A2(\converter/_111_ ),
    .ZN(\converter/_128_ ));
 INV_X1 \converter/_197_  (.A(net11),
    .ZN(\converter/_129_ ));
 NAND2_X1 \converter/_198_  (.A1(\converter/_112_ ),
    .A2(\converter/_129_ ),
    .ZN(\converter/_130_ ));
 NAND2_X1 \converter/_199_  (.A1(\converter/_130_ ),
    .A2(\converter/_109_ ),
    .ZN(\converter/_131_ ));
 NAND2_X1 \converter/_200_  (.A1(\converter/_131_ ),
    .A2(\converter/_108_ ),
    .ZN(\converter/_132_ ));
 INV_X1 \converter/_201_  (.A(\converter/_132_ ),
    .ZN(\converter/_133_ ));
 NAND2_X2 \converter/_202_  (.A1(\converter/_128_ ),
    .A2(\converter/_133_ ),
    .ZN(\converter/_134_ ));
 INV_X4 \converter/_203_  (.A(\converter/_134_ ),
    .ZN(\converter/_135_ ));
 NOR2_X2 \converter/_204_  (.A1(\converter/_127_ ),
    .A2(\converter/_110_ ),
    .ZN(\converter/_136_ ));
 NAND3_X1 \converter/_205_  (.A1(\converter/_126_ ),
    .A2(\converter/_135_ ),
    .A3(\converter/_136_ ),
    .ZN(\converter/_137_ ));
 NOR2_X1 \converter/_206_  (.A1(net8),
    .A2(net1),
    .ZN(\converter/_138_ ));
 INV_X1 \converter/_207_  (.A(\converter/_138_ ),
    .ZN(\converter/_139_ ));
 NAND2_X1 \converter/_208_  (.A1(\converter/_121_ ),
    .A2(\converter/_139_ ),
    .ZN(\converter/_140_ ));
 NAND2_X1 \converter/_209_  (.A1(\converter/_137_ ),
    .A2(\converter/_140_ ),
    .ZN(\converter/_141_ ));
 INV_X2 \converter/_210_  (.A(\converter/_141_ ),
    .ZN(\converter/_142_ ));
 OAI21_X2 \converter/_211_  (.A(\converter/_099_ ),
    .B1(\converter/_128_ ),
    .B2(\converter/_139_ ),
    .ZN(\converter/_143_ ));
 INV_X1 \converter/_212_  (.A(\converter/_143_ ),
    .ZN(\converter/_144_ ));
 NAND2_X2 \converter/_213_  (.A1(\converter/_142_ ),
    .A2(\converter/_144_ ),
    .ZN(\converter/_145_ ));
 TAPCELL_X1 PHY_18 ();
 TAPCELL_X1 PHY_17 ();
 NAND3_X1 \converter/_216_  (.A1(\converter/_117_ ),
    .A2(\converter/_134_ ),
    .A3(\converter/_124_ ),
    .ZN(\converter/_148_ ));
 NAND2_X1 \converter/_217_  (.A1(net262),
    .A2(\converter/_135_ ),
    .ZN(\converter/_149_ ));
 NAND2_X4 \converter/_218_  (.A1(\converter/_148_ ),
    .A2(\converter/_149_ ),
    .ZN(\converter/_150_ ));
 TAPCELL_X1 PHY_16 ();
 INV_X1 \converter/_220_  (.A(net1),
    .ZN(\converter/_152_ ));
 NAND2_X1 \converter/_221_  (.A1(net264),
    .A2(\converter/_152_ ),
    .ZN(\converter/_153_ ));
 NAND3_X1 \converter/_222_  (.A1(\converter/_117_ ),
    .A2(\converter/_124_ ),
    .A3(\converter/_122_ ),
    .ZN(\converter/_154_ ));
 NAND2_X1 \converter/_223_  (.A1(\converter/_153_ ),
    .A2(\converter/_154_ ),
    .ZN(\converter/_155_ ));
 NOR2_X1 \converter/_224_  (.A1(\converter/_150_ ),
    .A2(\converter/_155_ ),
    .ZN(\converter/_156_ ));
 NAND3_X1 \converter/_225_  (.A1(\converter/_135_ ),
    .A2(\converter/_117_ ),
    .A3(\converter/_124_ ),
    .ZN(\converter/_157_ ));
 INV_X1 \converter/_226_  (.A(\converter/_136_ ),
    .ZN(\converter/_158_ ));
 NAND2_X1 \converter/_227_  (.A1(\converter/_157_ ),
    .A2(\converter/_158_ ),
    .ZN(\converter/_159_ ));
 NAND2_X2 \converter/_228_  (.A1(\converter/_137_ ),
    .A2(\converter/_159_ ),
    .ZN(\converter/_160_ ));
 NAND2_X1 \converter/_229_  (.A1(\converter/_156_ ),
    .A2(\converter/_160_ ),
    .ZN(\converter/_000_ ));
 OAI22_X2 \converter/_230_  (.A1(\converter/_145_ ),
    .A2(\converter/_000_ ),
    .B1(\converter/_122_ ),
    .B2(\converter/_099_ ),
    .ZN(\operand_fp16_fp32[14] ));
 NAND2_X1 \converter/_231_  (.A1(\converter/_100_ ),
    .A2(net9),
    .ZN(\converter/_001_ ));
 INV_X4 \converter/_232_  (.A(\converter/_145_ ),
    .ZN(\converter/_002_ ));
 NAND2_X1 \converter/_233_  (.A1(\converter/_002_ ),
    .A2(\converter/_160_ ),
    .ZN(\converter/_003_ ));
 NAND2_X1 \converter/_234_  (.A1(\converter/_126_ ),
    .A2(net1),
    .ZN(\converter/_004_ ));
 NAND2_X1 \converter/_235_  (.A1(\converter/_150_ ),
    .A2(\converter/_004_ ),
    .ZN(\converter/_005_ ));
 NAND2_X1 \converter/_236_  (.A1(net262),
    .A2(net8),
    .ZN(\converter/_006_ ));
 NAND3_X1 \converter/_237_  (.A1(net269),
    .A2(\converter/_124_ ),
    .A3(net9),
    .ZN(\converter/_007_ ));
 NAND2_X1 \converter/_238_  (.A1(\converter/_006_ ),
    .A2(\converter/_007_ ),
    .ZN(\converter/_008_ ));
 OAI21_X1 \converter/_239_  (.A(\converter/_005_ ),
    .B1(\converter/_150_ ),
    .B2(\converter/_008_ ),
    .ZN(\converter/_009_ ));
 OAI21_X1 \converter/_240_  (.A(\converter/_001_ ),
    .B1(\converter/_003_ ),
    .B2(\converter/_009_ ),
    .ZN(\operand_fp16_fp32[15] ));
 NAND2_X1 \converter/_241_  (.A1(\converter/_100_ ),
    .A2(net10),
    .ZN(\converter/_010_ ));
 NAND2_X1 \converter/_242_  (.A1(net263),
    .A2(net9),
    .ZN(\converter/_011_ ));
 NAND3_X1 \converter/_243_  (.A1(net269),
    .A2(\converter/_124_ ),
    .A3(net10),
    .ZN(\converter/_012_ ));
 NAND2_X1 \converter/_244_  (.A1(\converter/_011_ ),
    .A2(\converter/_012_ ),
    .ZN(\converter/_013_ ));
 INV_X1 \converter/_245_  (.A(\converter/_013_ ),
    .ZN(\converter/_014_ ));
 NAND2_X1 \converter/_246_  (.A1(\converter/_125_ ),
    .A2(\converter/_134_ ),
    .ZN(\converter/_015_ ));
 NAND2_X2 \converter/_247_  (.A1(\converter/_157_ ),
    .A2(\converter/_015_ ),
    .ZN(\converter/_016_ ));
 NAND2_X1 \converter/_248_  (.A1(\converter/_014_ ),
    .A2(\converter/_016_ ),
    .ZN(\converter/_017_ ));
 NAND2_X1 \converter/_249_  (.A1(\converter/_150_ ),
    .A2(\converter/_155_ ),
    .ZN(\converter/_018_ ));
 NAND2_X1 \converter/_250_  (.A1(\converter/_017_ ),
    .A2(\converter/_018_ ),
    .ZN(\converter/_019_ ));
 OAI21_X1 \converter/_251_  (.A(\converter/_010_ ),
    .B1(\converter/_003_ ),
    .B2(\converter/_019_ ),
    .ZN(\operand_fp16_fp32[16] ));
 INV_X2 \converter/_252_  (.A(\converter/_160_ ),
    .ZN(\converter/_020_ ));
 OAI21_X1 \converter/_253_  (.A(\converter/_020_ ),
    .B1(\converter/_150_ ),
    .B2(\converter/_004_ ),
    .ZN(\converter/_021_ ));
 NAND2_X1 \converter/_254_  (.A1(net262),
    .A2(net10),
    .ZN(\converter/_022_ ));
 NAND3_X1 \converter/_255_  (.A1(net269),
    .A2(\converter/_124_ ),
    .A3(net11),
    .ZN(\converter/_023_ ));
 NAND2_X1 \converter/_256_  (.A1(\converter/_022_ ),
    .A2(\converter/_023_ ),
    .ZN(\converter/_024_ ));
 NAND2_X1 \converter/_257_  (.A1(\converter/_016_ ),
    .A2(\converter/_024_ ),
    .ZN(\converter/_025_ ));
 NAND2_X1 \converter/_258_  (.A1(\converter/_150_ ),
    .A2(\converter/_008_ ),
    .ZN(\converter/_026_ ));
 NAND3_X1 \converter/_259_  (.A1(\converter/_160_ ),
    .A2(\converter/_025_ ),
    .A3(\converter/_026_ ),
    .ZN(\converter/_027_ ));
 NAND3_X1 \converter/_260_  (.A1(\converter/_021_ ),
    .A2(\converter/_002_ ),
    .A3(\converter/_027_ ),
    .ZN(\converter/_028_ ));
 NAND2_X1 \converter/_261_  (.A1(\converter/_100_ ),
    .A2(net11),
    .ZN(\converter/_029_ ));
 NAND2_X1 \converter/_262_  (.A1(\converter/_028_ ),
    .A2(\converter/_029_ ),
    .ZN(\operand_fp16_fp32[17] ));
 NAND2_X1 \converter/_263_  (.A1(\converter/_100_ ),
    .A2(net12),
    .ZN(\converter/_030_ ));
 OR2_X1 \converter/_264_  (.A1(\converter/_156_ ),
    .A2(\converter/_160_ ),
    .ZN(\converter/_031_ ));
 NAND2_X1 \converter/_265_  (.A1(\converter/_031_ ),
    .A2(\converter/_002_ ),
    .ZN(\converter/_032_ ));
 NAND2_X1 \converter/_266_  (.A1(net263),
    .A2(net11),
    .ZN(\converter/_033_ ));
 NAND3_X1 \converter/_267_  (.A1(net270),
    .A2(\converter/_124_ ),
    .A3(net12),
    .ZN(\converter/_034_ ));
 NAND2_X1 \converter/_268_  (.A1(\converter/_033_ ),
    .A2(\converter/_034_ ),
    .ZN(\converter/_035_ ));
 NAND2_X1 \converter/_269_  (.A1(\converter/_016_ ),
    .A2(\converter/_035_ ),
    .ZN(\converter/_036_ ));
 NAND2_X1 \converter/_270_  (.A1(\converter/_150_ ),
    .A2(\converter/_013_ ),
    .ZN(\converter/_037_ ));
 NAND2_X1 \converter/_271_  (.A1(\converter/_036_ ),
    .A2(\converter/_037_ ),
    .ZN(\converter/_038_ ));
 NOR2_X1 \converter/_272_  (.A1(\converter/_038_ ),
    .A2(\converter/_020_ ),
    .ZN(\converter/_039_ ));
 OAI21_X2 \converter/_273_  (.A(\converter/_030_ ),
    .B1(\converter/_032_ ),
    .B2(\converter/_039_ ),
    .ZN(\operand_fp16_fp32[18] ));
 NAND2_X1 \converter/_274_  (.A1(net262),
    .A2(\converter/_112_ ),
    .ZN(\converter/_040_ ));
 INV_X1 \converter/_275_  (.A(net13),
    .ZN(\converter/_041_ ));
 NAND3_X1 \converter/_276_  (.A1(net269),
    .A2(\converter/_124_ ),
    .A3(\converter/_041_ ),
    .ZN(\converter/_042_ ));
 NAND2_X1 \converter/_277_  (.A1(\converter/_040_ ),
    .A2(\converter/_042_ ),
    .ZN(\converter/_043_ ));
 NAND2_X1 \converter/_278_  (.A1(\converter/_016_ ),
    .A2(\converter/_043_ ),
    .ZN(\converter/_044_ ));
 OAI21_X1 \converter/_279_  (.A(\converter/_044_ ),
    .B1(\converter/_016_ ),
    .B2(\converter/_024_ ),
    .ZN(\converter/_045_ ));
 NOR2_X1 \converter/_280_  (.A1(\converter/_045_ ),
    .A2(\converter/_145_ ),
    .ZN(\converter/_046_ ));
 NAND2_X1 \converter/_281_  (.A1(\converter/_009_ ),
    .A2(\converter/_020_ ),
    .ZN(\converter/_047_ ));
 NAND2_X1 \converter/_282_  (.A1(\converter/_046_ ),
    .A2(\converter/_047_ ),
    .ZN(\converter/_048_ ));
 NAND2_X1 \converter/_283_  (.A1(\converter/_100_ ),
    .A2(net13),
    .ZN(\converter/_049_ ));
 NAND2_X1 \converter/_284_  (.A1(\converter/_048_ ),
    .A2(\converter/_049_ ),
    .ZN(\operand_fp16_fp32[19] ));
 NAND2_X1 \converter/_285_  (.A1(\converter/_019_ ),
    .A2(\converter/_020_ ),
    .ZN(\converter/_050_ ));
 INV_X1 \converter/_286_  (.A(\converter/_035_ ),
    .ZN(\converter/_051_ ));
 NAND2_X1 \converter/_287_  (.A1(\converter/_051_ ),
    .A2(\converter/_150_ ),
    .ZN(\converter/_052_ ));
 NAND2_X1 \converter/_288_  (.A1(net262),
    .A2(\converter/_041_ ),
    .ZN(\converter/_053_ ));
 NAND3_X1 \converter/_289_  (.A1(net269),
    .A2(\converter/_124_ ),
    .A3(\converter/_105_ ),
    .ZN(\converter/_054_ ));
 NAND2_X1 \converter/_290_  (.A1(\converter/_053_ ),
    .A2(\converter/_054_ ),
    .ZN(\converter/_055_ ));
 NAND2_X1 \converter/_291_  (.A1(\converter/_016_ ),
    .A2(\converter/_055_ ),
    .ZN(\converter/_056_ ));
 NAND2_X1 \converter/_292_  (.A1(\converter/_052_ ),
    .A2(\converter/_056_ ),
    .ZN(\converter/_057_ ));
 NAND2_X1 \converter/_293_  (.A1(\converter/_057_ ),
    .A2(\converter/_160_ ),
    .ZN(\converter/_058_ ));
 NAND3_X1 \converter/_294_  (.A1(\converter/_050_ ),
    .A2(\converter/_058_ ),
    .A3(\converter/_099_ ),
    .ZN(\converter/_059_ ));
 NAND2_X1 \converter/_295_  (.A1(\converter/_100_ ),
    .A2(net14),
    .ZN(\converter/_060_ ));
 NAND2_X1 \converter/_296_  (.A1(\converter/_059_ ),
    .A2(\converter/_060_ ),
    .ZN(\operand_fp16_fp32[20] ));
 NAND2_X1 \converter/_297_  (.A1(net262),
    .A2(\converter/_105_ ),
    .ZN(\converter/_061_ ));
 INV_X1 \converter/_298_  (.A(net15),
    .ZN(\converter/_062_ ));
 NAND3_X1 \converter/_299_  (.A1(\converter/_117_ ),
    .A2(\converter/_124_ ),
    .A3(\converter/_062_ ),
    .ZN(\converter/_063_ ));
 NAND2_X1 \converter/_300_  (.A1(\converter/_061_ ),
    .A2(\converter/_063_ ),
    .ZN(\converter/_064_ ));
 NAND2_X1 \converter/_301_  (.A1(\converter/_016_ ),
    .A2(\converter/_064_ ),
    .ZN(\converter/_065_ ));
 NAND2_X1 \converter/_302_  (.A1(\converter/_150_ ),
    .A2(\converter/_043_ ),
    .ZN(\converter/_066_ ));
 NAND2_X1 \converter/_303_  (.A1(\converter/_065_ ),
    .A2(\converter/_066_ ),
    .ZN(\converter/_067_ ));
 NAND2_X1 \converter/_304_  (.A1(\converter/_067_ ),
    .A2(\converter/_142_ ),
    .ZN(\converter/_068_ ));
 INV_X1 \converter/_305_  (.A(\converter/_068_ ),
    .ZN(\converter/_069_ ));
 NAND2_X1 \converter/_306_  (.A1(\converter/_025_ ),
    .A2(\converter/_026_ ),
    .ZN(\converter/_070_ ));
 NAND2_X1 \converter/_307_  (.A1(\converter/_070_ ),
    .A2(\converter/_020_ ),
    .ZN(\converter/_071_ ));
 NAND2_X1 \converter/_308_  (.A1(\converter/_069_ ),
    .A2(\converter/_071_ ),
    .ZN(\converter/_072_ ));
 NAND4_X1 \converter/_309_  (.A1(\converter/_126_ ),
    .A2(net1),
    .A3(\converter/_135_ ),
    .A4(\converter/_136_ ),
    .ZN(\converter/_073_ ));
 AOI21_X1 \converter/_310_  (.A(\converter/_143_ ),
    .B1(\converter/_141_ ),
    .B2(\converter/_073_ ),
    .ZN(\converter/_074_ ));
 NAND2_X1 \converter/_311_  (.A1(\converter/_072_ ),
    .A2(\converter/_074_ ),
    .ZN(\converter/_075_ ));
 NAND2_X1 \converter/_312_  (.A1(\converter/_100_ ),
    .A2(net15),
    .ZN(\converter/_076_ ));
 NAND2_X1 \converter/_313_  (.A1(\converter/_075_ ),
    .A2(\converter/_076_ ),
    .ZN(\operand_fp16_fp32[21] ));
 NAND2_X1 \converter/_314_  (.A1(net262),
    .A2(net15),
    .ZN(\converter/_077_ ));
 NAND2_X1 \converter/_315_  (.A1(\converter/_016_ ),
    .A2(\converter/_077_ ),
    .ZN(\converter/_078_ ));
 NAND2_X1 \converter/_316_  (.A1(\converter/_150_ ),
    .A2(\converter/_055_ ),
    .ZN(\converter/_079_ ));
 NAND2_X1 \converter/_317_  (.A1(\converter/_078_ ),
    .A2(\converter/_079_ ),
    .ZN(\converter/_080_ ));
 NAND2_X1 \converter/_318_  (.A1(\converter/_080_ ),
    .A2(\converter/_142_ ),
    .ZN(\converter/_081_ ));
 INV_X1 \converter/_319_  (.A(\converter/_081_ ),
    .ZN(\converter/_082_ ));
 NAND2_X1 \converter/_320_  (.A1(\converter/_038_ ),
    .A2(\converter/_020_ ),
    .ZN(\converter/_083_ ));
 NAND2_X1 \converter/_321_  (.A1(\converter/_082_ ),
    .A2(\converter/_083_ ),
    .ZN(\converter/_084_ ));
 AOI21_X1 \converter/_322_  (.A(\converter/_143_ ),
    .B1(\converter/_000_ ),
    .B2(\converter/_141_ ),
    .ZN(\converter/_085_ ));
 NAND2_X1 \converter/_323_  (.A1(\converter/_084_ ),
    .A2(\converter/_085_ ),
    .ZN(\converter/_086_ ));
 NAND2_X1 \converter/_324_  (.A1(\converter/_100_ ),
    .A2(net16),
    .ZN(\converter/_087_ ));
 NAND2_X1 \converter/_325_  (.A1(\converter/_086_ ),
    .A2(\converter/_087_ ),
    .ZN(\operand_fp16_fp32[22] ));
 OAI21_X2 \converter/_326_  (.A(\converter/_096_ ),
    .B1(\converter/_100_ ),
    .B2(\converter/_125_ ),
    .ZN(\operand_fp16_fp32[23] ));
 OAI21_X2 \converter/_327_  (.A(\converter/_095_ ),
    .B1(\converter/_016_ ),
    .B2(\converter/_100_ ),
    .ZN(\operand_fp16_fp32[24] ));
 NAND2_X1 \converter/_328_  (.A1(\converter/_015_ ),
    .A2(\converter/_136_ ),
    .ZN(\converter/_088_ ));
 NAND3_X1 \converter/_329_  (.A1(\converter/_125_ ),
    .A2(\converter/_134_ ),
    .A3(\converter/_158_ ),
    .ZN(\converter/_089_ ));
 NAND3_X1 \converter/_330_  (.A1(\converter/_088_ ),
    .A2(\converter/_089_ ),
    .A3(\converter/_099_ ),
    .ZN(\converter/_090_ ));
 INV_X1 \converter/_331_  (.A(net4),
    .ZN(\converter/_091_ ));
 NAND2_X1 \converter/_332_  (.A1(\converter/_090_ ),
    .A2(\converter/_091_ ),
    .ZN(\operand_fp16_fp32[25] ));
 INV_X1 \converter/_333_  (.A(net5),
    .ZN(\converter/_092_ ));
 XOR2_X1 \converter/_334_  (.A(\converter/_089_ ),
    .B(\converter/_140_ ),
    .Z(\converter/_093_ ));
 OAI21_X2 \converter/_335_  (.A(\converter/_092_ ),
    .B1(\converter/_093_ ),
    .B2(\converter/_100_ ),
    .ZN(\operand_fp16_fp32[26] ));
 NAND2_X1 \converter/_336_  (.A1(\converter/_099_ ),
    .A2(net16),
    .ZN(\converter/_094_ ));
 OAI21_X1 \converter/_337_  (.A(\converter/_094_ ),
    .B1(net6),
    .B2(\converter/_099_ ),
    .ZN(\operand_fp16_fp32[27] ));
 OAI21_X2 \converter/_338_  (.A(\converter/_143_ ),
    .B1(net6),
    .B2(\converter/_099_ ),
    .ZN(\operand_fp16_fp32[29] ));
 TAPCELL_X1 PHY_15 ();
 BUF_X8 split1 (.A(net242),
    .Z(net239));
 TAPCELL_X1 PHY_14 ();
 TAPCELL_X1 PHY_13 ();
 TAPCELL_X1 PHY_12 ();
 TAPCELL_X1 PHY_11 ();
 TAPCELL_X1 PHY_10 ();
 TAPCELL_X1 PHY_9 ();
 TAPCELL_X1 PHY_8 ();
 TAPCELL_X1 PHY_7 ();
 TAPCELL_X1 PHY_6 ();
 TAPCELL_X1 PHY_5 ();
 TAPCELL_X1 PHY_4 ();
 TAPCELL_X1 PHY_3 ();
 TAPCELL_X1 PHY_2 ();
 TAPCELL_X1 PHY_1 ();
 TAPCELL_X1 PHY_0 ();
 LOGIC0_X1 \adder/norm/LOD/_217__86  (.Z(net86));
 LOGIC0_X1 \adder/norm/LOD/_218__87  (.Z(net87));
 LOGIC0_X1 \adder/norm/LOD/_218__88  (.Z(net88));
 LOGIC0_X1 \adder/norm/LOD/_228__89  (.Z(net89));
 LOGIC0_X1 \adder/norm/LOD/_228__90  (.Z(net90));
 LOGIC0_X1 \adder/norm/LOD/_229__91  (.Z(net91));
 LOGIC0_X1 \adder/norm/LOD/_230__92  (.Z(net92));
 LOGIC0_X1 \adder/norm/LOD/_239__93  (.Z(net93));
 LOGIC0_X1 \adder/norm/LOD/_239__94  (.Z(net94));
 LOGIC0_X1 \adder/norm/LOD/_240__95  (.Z(net95));
 LOGIC0_X1 \adder/norm/LOD/_241__96  (.Z(net96));
 LOGIC0_X1 \adder/norm/LOD/_243__97  (.Z(net97));
 LOGIC0_X1 \adder/norm/LOD/_243__98  (.Z(net98));
 LOGIC0_X1 \adder/norm/LOD/_245__99  (.Z(net99));
 LOGIC0_X1 \adder/norm/LOD/_246__100  (.Z(net100));
 LOGIC0_X1 \adder/norm/LOD/_247__101  (.Z(net101));
 LOGIC0_X1 \adder/norm/LOD/_249__102  (.Z(net102));
 LOGIC0_X1 \adder/norm/LOD/_249__103  (.Z(net103));
 LOGIC0_X1 \adder/norm/LOD/_250__104  (.Z(net104));
 LOGIC0_X1 \adder/norm/LOD/_255__105  (.Z(net105));
 LOGIC0_X1 \adder/norm/LOD/_255__106  (.Z(net106));
 LOGIC0_X1 \adder/norm/LOD/_256__107  (.Z(net107));
 LOGIC0_X1 \adder/norm/LOD/_257__108  (.Z(net108));
 LOGIC0_X1 \adder/norm/LOD/_259__109  (.Z(net109));
 LOGIC0_X1 \adder/norm/LOD/_260__110  (.Z(net110));
 LOGIC0_X1 \adder/norm/LOD/_260__111  (.Z(net111));
 LOGIC0_X1 \adder/norm/LOD/_262__112  (.Z(net112));
 LOGIC0_X1 \adder/norm/LOD/_263__113  (.Z(net113));
 LOGIC0_X1 \adder/norm/LOD/_264__114  (.Z(net114));
 LOGIC0_X1 \adder/norm/LOD/_269__115  (.Z(net115));
 LOGIC0_X1 \adder/norm/LOD/_269__116  (.Z(net116));
 LOGIC0_X1 \adder/norm/LOD/_270__117  (.Z(net117));
 LOGIC0_X1 \adder/norm/LOD/_270__118  (.Z(net118));
 LOGIC0_X1 \adder/norm/LOD/_299__119  (.Z(net119));
 LOGIC0_X1 \adder/norm/LOD/_299__120  (.Z(net120));
 LOGIC0_X1 \adder/norm/_1529__121  (.Z(net121));
 LOGIC0_X1 \adder/norm/_1531__122  (.Z(net122));
 LOGIC0_X1 \adder/norm/_1533__123  (.Z(net123));
 LOGIC0_X1 \adder/norm/_1551__124  (.Z(net124));
 LOGIC0_X1 \adder/norm/_1634__125  (.Z(net125));
 LOGIC0_X1 \adder/norm/_1635__126  (.Z(net126));
 LOGIC0_X1 \adder/norm/_1669__127  (.Z(net127));
 LOGIC0_X1 \adder/norm/_1674__128  (.Z(net128));
 LOGIC0_X1 \adder/norm/_1679__129  (.Z(net129));
 LOGIC0_X1 \adder/norm/_1681__130  (.Z(net130));
 LOGIC0_X1 \adder/norm/_1688__131  (.Z(net131));
 LOGIC0_X1 \adder/norm/_1690__132  (.Z(net132));
 LOGIC0_X1 \adder/norm/_1694__133  (.Z(net133));
 LOGIC0_X1 \adder/norm/_1696__134  (.Z(net134));
 LOGIC0_X1 \adder/norm/_1701__135  (.Z(net135));
 LOGIC0_X1 \adder/norm/_1703__136  (.Z(net136));
 LOGIC0_X1 \adder/norm/_1707__137  (.Z(net137));
 LOGIC0_X1 \adder/norm/_1710__138  (.Z(net138));
 LOGIC0_X1 \adder/norm/_1713__139  (.Z(net139));
 LOGIC0_X1 \adder/norm/_1715__140  (.Z(net140));
 LOGIC0_X1 \adder/norm/_1719__141  (.Z(net141));
 LOGIC0_X1 \adder/norm/_1720__142  (.Z(net142));
 LOGIC0_X1 \adder/norm/_1782__143  (.Z(net143));
 LOGIC0_X1 \adder/norm/_1785__144  (.Z(net144));
 LOGIC0_X1 \adder/norm/_1814__145  (.Z(net145));
 LOGIC0_X1 \adder/norm/_1816__146  (.Z(net146));
 LOGIC0_X1 \adder/norm/_1817__147  (.Z(net147));
 LOGIC0_X1 \adder/norm/_1846__148  (.Z(net148));
 LOGIC0_X1 \adder/norm/_1847__149  (.Z(net149));
 LOGIC0_X1 \adder/norm/_1850__150  (.Z(net150));
 LOGIC0_X1 \adder/norm/_1851__151  (.Z(net151));
 LOGIC0_X1 \adder/norm/_1853__152  (.Z(net152));
 LOGIC0_X1 \adder/norm/_1854__153  (.Z(net153));
 LOGIC0_X1 \adder/norm/_1858__154  (.Z(net154));
 LOGIC0_X1 \adder/norm/_1859__155  (.Z(net155));
 LOGIC0_X1 \adder/norm/_1861__156  (.Z(net156));
 LOGIC0_X1 \adder/norm/_1862__157  (.Z(net157));
 LOGIC0_X1 \adder/norm/_1866__158  (.Z(net158));
 LOGIC0_X1 \adder/norm/_1867__159  (.Z(net159));
 LOGIC0_X1 \adder/norm/_1869__160  (.Z(net160));
 LOGIC0_X1 \adder/norm/_1870__161  (.Z(net161));
 LOGIC0_X1 \adder/norm/_1912__162  (.Z(net162));
 LOGIC0_X1 \adder/norm/_2002__163  (.Z(net163));
 LOGIC0_X1 \adder/norm/_2004__164  (.Z(net164));
 LOGIC0_X1 \adder/norm/_2489__165  (.Z(net165));
 LOGIC0_X1 \adder/norm/_2536__166  (.Z(net166));
 LOGIC0_X1 \adder/norm/_2626__167  (.Z(net167));
 LOGIC0_X1 \adder/norm/_2630__168  (.Z(net168));
 LOGIC0_X1 \adder/norm/_2635__169  (.Z(net169));
 LOGIC0_X1 \adder/norm/_2637__170  (.Z(net170));
 LOGIC0_X1 \adder/norm/_2751__171  (.Z(net171));
 LOGIC0_X1 \adder/norm/_2756__172  (.Z(net172));
 LOGIC0_X1 \adder/norm/_2758__173  (.Z(net173));
 LOGIC0_X1 \adder/norm/_2764__174  (.Z(net174));
 LOGIC0_X1 \adder/norm/_2767__175  (.Z(net175));
 LOGIC0_X1 \adder/norm/_2768__176  (.Z(net176));
 LOGIC0_X1 \adder/norm/_2772__177  (.Z(net177));
 LOGIC0_X1 \adder/norm/_2774__178  (.Z(net178));
 LOGIC0_X1 \adder/norm/_2782__179  (.Z(net179));
 LOGIC0_X1 \adder/norm/_2798__180  (.Z(net180));
 LOGIC0_X1 \adder/norm/_2801__181  (.Z(net181));
 LOGIC0_X1 \adder/norm/_2894__182  (.Z(net182));
 LOGIC0_X1 \adder/norm/_2894__183  (.Z(net183));
 LOGIC0_X1 \adder/norm/_2894__184  (.Z(net184));
 LOGIC0_X1 \adder/norm/_2894__185  (.Z(net185));
 LOGIC0_X1 \adder/norm/_2895__186  (.Z(net186));
 LOGIC0_X1 \adder/norm/_2895__187  (.Z(net187));
 LOGIC0_X1 \adder/norm/_2895__188  (.Z(net188));
 LOGIC0_X1 \adder/norm/_2895__189  (.Z(net189));
 LOGIC0_X1 \adder/norm/_2896__190  (.Z(net190));
 LOGIC0_X1 \adder/norm/_2896__191  (.Z(net191));
 LOGIC0_X1 \adder/norm/_2896__192  (.Z(net192));
 LOGIC0_X1 \adder/norm/_2896__193  (.Z(net193));
 LOGIC0_X1 \adder/norm/_2897__194  (.Z(net194));
 LOGIC0_X1 \adder/norm/_2897__195  (.Z(net195));
 LOGIC0_X1 \adder/norm/_2897__196  (.Z(net196));
 LOGIC0_X1 \adder/norm/_2897__197  (.Z(net197));
 LOGIC0_X1 \adder/norm/_2899__198  (.Z(net198));
 LOGIC0_X1 \adder/norm/_2899__199  (.Z(net199));
 LOGIC0_X1 \adder/norm/_2899__200  (.Z(net200));
 LOGIC0_X1 \adder/norm/_2899__201  (.Z(net201));
 LOGIC0_X1 \adder/adder/_1356__203  (.Z(net203));
 LOGIC0_X1 \adder/adder/_1477__204  (.Z(net204));
 LOGIC0_X1 \adder/adder/_1492__205  (.Z(net205));
 LOGIC0_X1 \adder/adder/_1513__206  (.Z(net206));
 LOGIC0_X1 \adder/adder/_1789__207  (.Z(net207));
 LOGIC0_X1 \adder/adder/_1804__208  (.Z(net208));
 LOGIC0_X1 \adder/adder/_1837__209  (.Z(net209));
 LOGIC0_X1 \adder/adder/_1857__210  (.Z(net210));
 LOGIC0_X1 \adder/adder/_1888__211  (.Z(net211));
 LOGIC0_X1 \adder/adder/_1898__212  (.Z(net212));
 LOGIC0_X1 \adder/adder/_1921__213  (.Z(net213));
 LOGIC0_X1 \adder/adder/_1931__214  (.Z(net214));
 LOGIC0_X1 \adder/adder/_1939__215  (.Z(net215));
 LOGIC0_X1 \adder/adder/_1948__216  (.Z(net216));
 LOGIC0_X1 \adder/adder/_2164__217  (.Z(net217));
 LOGIC0_X1 \adder/adder/_2167__218  (.Z(net218));
 LOGIC0_X1 \adder/adder/_2168__219  (.Z(net219));
 LOGIC0_X1 \adder/adder/_2171__220  (.Z(net220));
 LOGIC0_X1 \adder/adder/_2172__221  (.Z(net221));
 LOGIC0_X1 \adder/adder/_2173__222  (.Z(net222));
 LOGIC0_X1 \adder/adder/_2176__223  (.Z(net223));
 LOGIC0_X1 \adder/adder/_2177__224  (.Z(net224));
 LOGIC0_X1 \adder/adder/_2181__225  (.Z(net225));
 LOGIC0_X1 \adder/adder/_2184__226  (.Z(net226));
 LOGIC0_X1 \adder/adder/_2186__227  (.Z(net227));
 LOGIC0_X1 \adder/adder/_2188__228  (.Z(net228));
 LOGIC0_X1 \adder/adder/_2191__229  (.Z(net229));
 LOGIC0_X1 \adder/adder/_2205__230  (.Z(net230));
 LOGIC0_X1 \adder/adder/_2211__231  (.Z(net231));
 LOGIC0_X1 \adder/adder/_2212__232  (.Z(net232));
 LOGIC0_X1 \adder/adder/_2214__233  (.Z(net233));
 LOGIC0_X1 \adder/adder/_2217__234  (.Z(net234));
 LOGIC0_X1 \adder/adder/_2219__235  (.Z(net235));
 LOGIC0_X1 \adder/adder/_2220__236  (.Z(net236));
 LOGIC0_X1 \adder/adder/_2223__237  (.Z(net237));
 LOGIC0_X1 \adder/adder/_2238__238  (.Z(net238));
 BUF_X8 split2 (.A(net241),
    .Z(net240));
 BUF_X8 split3 (.A(\adder/norm/_0638_ ),
    .Z(net241));
 BUF_X8 split4 (.A(net251),
    .Z(net242));
 CLKBUF_X3 split5 (.A(\adder/norm/_0638_ ),
    .Z(net243));
 BUF_X4 split6 (.A(\adder/norm/_0658_ ),
    .Z(net244));
 BUF_X4 split7 (.A(net251),
    .Z(net245));
 CLKBUF_X3 split8 (.A(\adder/norm/_0638_ ),
    .Z(net246));
 CLKBUF_X3 split9 (.A(net256),
    .Z(net247));
 BUF_X4 split10 (.A(\adder/norm/_0082_ ),
    .Z(net248));
 CLKBUF_X3 split11 (.A(\adder/norm/_0658_ ),
    .Z(net249));
 BUF_X8 split12 (.A(\adder/norm/_0717_ ),
    .Z(net250));
 CLKBUF_X3 split13 (.A(\adder/adder/_0413_ ),
    .Z(net251));
 CLKBUF_X3 split14 (.A(\adder/adder/_0420_ ),
    .Z(net252));
 CLKBUF_X3 split15 (.A(\adder/adder/_0443_ ),
    .Z(net253));
 BUF_X4 split16 (.A(\adder/adder/_0458_ ),
    .Z(net254));
 BUF_X4 split17 (.A(\adder/adder/_0506_ ),
    .Z(net255));
 BUF_X4 split18 (.A(\adder/norm/_0659_ ),
    .Z(net256));
 BUF_X4 split19 (.A(\adder/norm/_0622_ ),
    .Z(net257));
 CLKBUF_X2 rebuffer20 (.A(\adder/norm/_0670_ ),
    .Z(net258));
 BUF_X8 rebuffer21 (.A(\adder/norm/_0638_ ),
    .Z(net259));
 BUF_X4 split22 (.A(\adder/norm/_0082_ ),
    .Z(net260));
 BUF_X4 rebuffer23 (.A(\adder/norm/_0082_ ),
    .Z(net261));
 CLKBUF_X3 rebuffer24 (.A(\converter/_125_ ),
    .Z(net262));
 CLKBUF_X1 rebuffer25 (.A(net262),
    .Z(net263));
 CLKBUF_X1 rebuffer26 (.A(net262),
    .Z(net264));
 BUF_X2 rebuffer27 (.A(\adder/adder/_0420_ ),
    .Z(net265));
 CLKBUF_X2 rebuffer28 (.A(\adder/adder/_0443_ ),
    .Z(net266));
 CLKBUF_X3 split29 (.A(\adder/adder/_0449_ ),
    .Z(net267));
 BUF_X2 split30 (.A(\adder/norm/_0658_ ),
    .Z(net268));
 CLKBUF_X1 rebuffer31 (.A(\converter/_117_ ),
    .Z(net269));
 CLKBUF_X1 rebuffer32 (.A(net269),
    .Z(net270));
 BUF_X4 split33 (.A(net84),
    .Z(net271));
 BUF_X2 split34 (.A(\adder/adder/_0458_ ),
    .Z(net272));
 FILLCELL_X32 FILLER_0_0_1 ();
 FILLCELL_X32 FILLER_0_0_33 ();
 FILLCELL_X32 FILLER_0_0_65 ();
 FILLCELL_X32 FILLER_0_0_97 ();
 FILLCELL_X8 FILLER_0_0_129 ();
 FILLCELL_X4 FILLER_0_0_137 ();
 FILLCELL_X4 FILLER_0_0_144 ();
 FILLCELL_X1 FILLER_0_0_148 ();
 FILLCELL_X8 FILLER_0_0_155 ();
 FILLCELL_X4 FILLER_0_0_163 ();
 FILLCELL_X1 FILLER_0_0_167 ();
 FILLCELL_X4 FILLER_0_0_171 ();
 FILLCELL_X1 FILLER_0_0_175 ();
 FILLCELL_X1 FILLER_0_0_179 ();
 FILLCELL_X4 FILLER_0_0_192 ();
 FILLCELL_X2 FILLER_0_0_196 ();
 FILLCELL_X4 FILLER_0_0_201 ();
 FILLCELL_X2 FILLER_0_0_205 ();
 FILLCELL_X1 FILLER_0_0_207 ();
 FILLCELL_X32 FILLER_0_0_211 ();
 FILLCELL_X32 FILLER_0_0_243 ();
 FILLCELL_X32 FILLER_0_0_275 ();
 FILLCELL_X32 FILLER_0_0_307 ();
 FILLCELL_X32 FILLER_0_0_339 ();
 FILLCELL_X32 FILLER_0_0_371 ();
 FILLCELL_X32 FILLER_0_0_403 ();
 FILLCELL_X32 FILLER_0_0_435 ();
 FILLCELL_X1 FILLER_0_0_467 ();
 FILLCELL_X32 FILLER_0_1_1 ();
 FILLCELL_X32 FILLER_0_1_33 ();
 FILLCELL_X32 FILLER_0_1_65 ();
 FILLCELL_X32 FILLER_0_1_97 ();
 FILLCELL_X32 FILLER_0_1_129 ();
 FILLCELL_X32 FILLER_0_1_161 ();
 FILLCELL_X16 FILLER_0_1_193 ();
 FILLCELL_X32 FILLER_0_1_212 ();
 FILLCELL_X32 FILLER_0_1_244 ();
 FILLCELL_X32 FILLER_0_1_276 ();
 FILLCELL_X32 FILLER_0_1_308 ();
 FILLCELL_X32 FILLER_0_1_340 ();
 FILLCELL_X32 FILLER_0_1_372 ();
 FILLCELL_X32 FILLER_0_1_404 ();
 FILLCELL_X32 FILLER_0_1_436 ();
 FILLCELL_X32 FILLER_0_2_1 ();
 FILLCELL_X32 FILLER_0_2_33 ();
 FILLCELL_X32 FILLER_0_2_65 ();
 FILLCELL_X32 FILLER_0_2_97 ();
 FILLCELL_X32 FILLER_0_2_129 ();
 FILLCELL_X32 FILLER_0_2_161 ();
 FILLCELL_X32 FILLER_0_2_193 ();
 FILLCELL_X32 FILLER_0_2_225 ();
 FILLCELL_X32 FILLER_0_2_257 ();
 FILLCELL_X32 FILLER_0_2_289 ();
 FILLCELL_X32 FILLER_0_2_321 ();
 FILLCELL_X32 FILLER_0_2_353 ();
 FILLCELL_X32 FILLER_0_2_385 ();
 FILLCELL_X32 FILLER_0_2_417 ();
 FILLCELL_X16 FILLER_0_2_449 ();
 FILLCELL_X2 FILLER_0_2_465 ();
 FILLCELL_X1 FILLER_0_2_467 ();
 FILLCELL_X32 FILLER_0_3_1 ();
 FILLCELL_X32 FILLER_0_3_33 ();
 FILLCELL_X32 FILLER_0_3_65 ();
 FILLCELL_X32 FILLER_0_3_97 ();
 FILLCELL_X32 FILLER_0_3_129 ();
 FILLCELL_X32 FILLER_0_3_161 ();
 FILLCELL_X32 FILLER_0_3_193 ();
 FILLCELL_X32 FILLER_0_3_225 ();
 FILLCELL_X32 FILLER_0_3_257 ();
 FILLCELL_X32 FILLER_0_3_289 ();
 FILLCELL_X32 FILLER_0_3_321 ();
 FILLCELL_X32 FILLER_0_3_353 ();
 FILLCELL_X32 FILLER_0_3_385 ();
 FILLCELL_X32 FILLER_0_3_417 ();
 FILLCELL_X16 FILLER_0_3_449 ();
 FILLCELL_X2 FILLER_0_3_465 ();
 FILLCELL_X1 FILLER_0_3_467 ();
 FILLCELL_X32 FILLER_0_4_1 ();
 FILLCELL_X32 FILLER_0_4_33 ();
 FILLCELL_X32 FILLER_0_4_65 ();
 FILLCELL_X32 FILLER_0_4_97 ();
 FILLCELL_X32 FILLER_0_4_129 ();
 FILLCELL_X32 FILLER_0_4_161 ();
 FILLCELL_X32 FILLER_0_4_193 ();
 FILLCELL_X32 FILLER_0_4_225 ();
 FILLCELL_X32 FILLER_0_4_257 ();
 FILLCELL_X32 FILLER_0_4_289 ();
 FILLCELL_X32 FILLER_0_4_321 ();
 FILLCELL_X32 FILLER_0_4_353 ();
 FILLCELL_X32 FILLER_0_4_385 ();
 FILLCELL_X32 FILLER_0_4_417 ();
 FILLCELL_X16 FILLER_0_4_449 ();
 FILLCELL_X2 FILLER_0_4_465 ();
 FILLCELL_X1 FILLER_0_4_467 ();
 FILLCELL_X32 FILLER_0_5_1 ();
 FILLCELL_X32 FILLER_0_5_33 ();
 FILLCELL_X32 FILLER_0_5_65 ();
 FILLCELL_X32 FILLER_0_5_97 ();
 FILLCELL_X32 FILLER_0_5_129 ();
 FILLCELL_X8 FILLER_0_5_161 ();
 FILLCELL_X1 FILLER_0_5_169 ();
 FILLCELL_X32 FILLER_0_5_172 ();
 FILLCELL_X32 FILLER_0_5_204 ();
 FILLCELL_X32 FILLER_0_5_236 ();
 FILLCELL_X32 FILLER_0_5_268 ();
 FILLCELL_X32 FILLER_0_5_300 ();
 FILLCELL_X32 FILLER_0_5_332 ();
 FILLCELL_X32 FILLER_0_5_364 ();
 FILLCELL_X32 FILLER_0_5_396 ();
 FILLCELL_X32 FILLER_0_5_428 ();
 FILLCELL_X8 FILLER_0_5_460 ();
 FILLCELL_X32 FILLER_0_6_1 ();
 FILLCELL_X32 FILLER_0_6_33 ();
 FILLCELL_X32 FILLER_0_6_65 ();
 FILLCELL_X32 FILLER_0_6_97 ();
 FILLCELL_X32 FILLER_0_6_129 ();
 FILLCELL_X16 FILLER_0_6_161 ();
 FILLCELL_X4 FILLER_0_6_177 ();
 FILLCELL_X1 FILLER_0_6_181 ();
 FILLCELL_X32 FILLER_0_6_184 ();
 FILLCELL_X32 FILLER_0_6_216 ();
 FILLCELL_X32 FILLER_0_6_248 ();
 FILLCELL_X32 FILLER_0_6_280 ();
 FILLCELL_X32 FILLER_0_6_312 ();
 FILLCELL_X32 FILLER_0_6_344 ();
 FILLCELL_X32 FILLER_0_6_376 ();
 FILLCELL_X32 FILLER_0_6_408 ();
 FILLCELL_X16 FILLER_0_6_440 ();
 FILLCELL_X8 FILLER_0_6_456 ();
 FILLCELL_X4 FILLER_0_6_464 ();
 FILLCELL_X32 FILLER_0_7_1 ();
 FILLCELL_X32 FILLER_0_7_33 ();
 FILLCELL_X32 FILLER_0_7_65 ();
 FILLCELL_X32 FILLER_0_7_97 ();
 FILLCELL_X4 FILLER_0_7_129 ();
 FILLCELL_X8 FILLER_0_7_145 ();
 FILLCELL_X2 FILLER_0_7_161 ();
 FILLCELL_X1 FILLER_0_7_163 ();
 FILLCELL_X16 FILLER_0_7_166 ();
 FILLCELL_X4 FILLER_0_7_182 ();
 FILLCELL_X32 FILLER_0_7_191 ();
 FILLCELL_X32 FILLER_0_7_223 ();
 FILLCELL_X32 FILLER_0_7_255 ();
 FILLCELL_X32 FILLER_0_7_287 ();
 FILLCELL_X32 FILLER_0_7_319 ();
 FILLCELL_X32 FILLER_0_7_351 ();
 FILLCELL_X32 FILLER_0_7_383 ();
 FILLCELL_X32 FILLER_0_7_415 ();
 FILLCELL_X16 FILLER_0_7_447 ();
 FILLCELL_X4 FILLER_0_7_463 ();
 FILLCELL_X1 FILLER_0_7_467 ();
 FILLCELL_X32 FILLER_0_8_1 ();
 FILLCELL_X32 FILLER_0_8_33 ();
 FILLCELL_X32 FILLER_0_8_65 ();
 FILLCELL_X8 FILLER_0_8_97 ();
 FILLCELL_X1 FILLER_0_8_105 ();
 FILLCELL_X1 FILLER_0_8_119 ();
 FILLCELL_X1 FILLER_0_8_167 ();
 FILLCELL_X2 FILLER_0_8_185 ();
 FILLCELL_X2 FILLER_0_8_196 ();
 FILLCELL_X1 FILLER_0_8_198 ();
 FILLCELL_X32 FILLER_0_8_203 ();
 FILLCELL_X32 FILLER_0_8_235 ();
 FILLCELL_X32 FILLER_0_8_267 ();
 FILLCELL_X32 FILLER_0_8_299 ();
 FILLCELL_X32 FILLER_0_8_331 ();
 FILLCELL_X32 FILLER_0_8_363 ();
 FILLCELL_X32 FILLER_0_8_395 ();
 FILLCELL_X32 FILLER_0_8_427 ();
 FILLCELL_X8 FILLER_0_8_459 ();
 FILLCELL_X1 FILLER_0_8_467 ();
 FILLCELL_X32 FILLER_0_9_1 ();
 FILLCELL_X32 FILLER_0_9_33 ();
 FILLCELL_X16 FILLER_0_9_65 ();
 FILLCELL_X4 FILLER_0_9_81 ();
 FILLCELL_X2 FILLER_0_9_85 ();
 FILLCELL_X16 FILLER_0_9_89 ();
 FILLCELL_X2 FILLER_0_9_105 ();
 FILLCELL_X8 FILLER_0_9_111 ();
 FILLCELL_X4 FILLER_0_9_119 ();
 FILLCELL_X8 FILLER_0_9_125 ();
 FILLCELL_X1 FILLER_0_9_133 ();
 FILLCELL_X2 FILLER_0_9_139 ();
 FILLCELL_X1 FILLER_0_9_141 ();
 FILLCELL_X4 FILLER_0_9_144 ();
 FILLCELL_X2 FILLER_0_9_150 ();
 FILLCELL_X1 FILLER_0_9_159 ();
 FILLCELL_X4 FILLER_0_9_162 ();
 FILLCELL_X8 FILLER_0_9_169 ();
 FILLCELL_X2 FILLER_0_9_177 ();
 FILLCELL_X1 FILLER_0_9_183 ();
 FILLCELL_X1 FILLER_0_9_186 ();
 FILLCELL_X32 FILLER_0_9_214 ();
 FILLCELL_X32 FILLER_0_9_246 ();
 FILLCELL_X32 FILLER_0_9_278 ();
 FILLCELL_X32 FILLER_0_9_310 ();
 FILLCELL_X32 FILLER_0_9_342 ();
 FILLCELL_X32 FILLER_0_9_374 ();
 FILLCELL_X32 FILLER_0_9_406 ();
 FILLCELL_X16 FILLER_0_9_438 ();
 FILLCELL_X8 FILLER_0_9_454 ();
 FILLCELL_X4 FILLER_0_9_462 ();
 FILLCELL_X2 FILLER_0_9_466 ();
 FILLCELL_X32 FILLER_0_10_1 ();
 FILLCELL_X16 FILLER_0_10_33 ();
 FILLCELL_X4 FILLER_0_10_49 ();
 FILLCELL_X2 FILLER_0_10_53 ();
 FILLCELL_X1 FILLER_0_10_55 ();
 FILLCELL_X4 FILLER_0_10_59 ();
 FILLCELL_X2 FILLER_0_10_92 ();
 FILLCELL_X1 FILLER_0_10_110 ();
 FILLCELL_X1 FILLER_0_10_114 ();
 FILLCELL_X2 FILLER_0_10_117 ();
 FILLCELL_X1 FILLER_0_10_122 ();
 FILLCELL_X8 FILLER_0_10_126 ();
 FILLCELL_X2 FILLER_0_10_140 ();
 FILLCELL_X4 FILLER_0_10_151 ();
 FILLCELL_X2 FILLER_0_10_155 ();
 FILLCELL_X1 FILLER_0_10_161 ();
 FILLCELL_X2 FILLER_0_10_164 ();
 FILLCELL_X2 FILLER_0_10_188 ();
 FILLCELL_X4 FILLER_0_10_216 ();
 FILLCELL_X32 FILLER_0_10_226 ();
 FILLCELL_X32 FILLER_0_10_258 ();
 FILLCELL_X32 FILLER_0_10_290 ();
 FILLCELL_X32 FILLER_0_10_322 ();
 FILLCELL_X32 FILLER_0_10_354 ();
 FILLCELL_X32 FILLER_0_10_386 ();
 FILLCELL_X32 FILLER_0_10_418 ();
 FILLCELL_X16 FILLER_0_10_450 ();
 FILLCELL_X2 FILLER_0_10_466 ();
 FILLCELL_X32 FILLER_0_11_1 ();
 FILLCELL_X2 FILLER_0_11_33 ();
 FILLCELL_X1 FILLER_0_11_35 ();
 FILLCELL_X1 FILLER_0_11_40 ();
 FILLCELL_X1 FILLER_0_11_47 ();
 FILLCELL_X8 FILLER_0_11_60 ();
 FILLCELL_X1 FILLER_0_11_68 ();
 FILLCELL_X1 FILLER_0_11_78 ();
 FILLCELL_X1 FILLER_0_11_93 ();
 FILLCELL_X4 FILLER_0_11_99 ();
 FILLCELL_X2 FILLER_0_11_103 ();
 FILLCELL_X1 FILLER_0_11_107 ();
 FILLCELL_X2 FILLER_0_11_121 ();
 FILLCELL_X1 FILLER_0_11_129 ();
 FILLCELL_X1 FILLER_0_11_149 ();
 FILLCELL_X2 FILLER_0_11_155 ();
 FILLCELL_X16 FILLER_0_11_163 ();
 FILLCELL_X4 FILLER_0_11_179 ();
 FILLCELL_X1 FILLER_0_11_190 ();
 FILLCELL_X2 FILLER_0_11_193 ();
 FILLCELL_X1 FILLER_0_11_199 ();
 FILLCELL_X32 FILLER_0_11_224 ();
 FILLCELL_X32 FILLER_0_11_256 ();
 FILLCELL_X32 FILLER_0_11_288 ();
 FILLCELL_X32 FILLER_0_11_320 ();
 FILLCELL_X32 FILLER_0_11_352 ();
 FILLCELL_X32 FILLER_0_11_384 ();
 FILLCELL_X32 FILLER_0_11_416 ();
 FILLCELL_X16 FILLER_0_11_448 ();
 FILLCELL_X4 FILLER_0_11_464 ();
 FILLCELL_X32 FILLER_0_12_1 ();
 FILLCELL_X2 FILLER_0_12_33 ();
 FILLCELL_X2 FILLER_0_12_38 ();
 FILLCELL_X2 FILLER_0_12_43 ();
 FILLCELL_X2 FILLER_0_12_48 ();
 FILLCELL_X1 FILLER_0_12_50 ();
 FILLCELL_X4 FILLER_0_12_54 ();
 FILLCELL_X1 FILLER_0_12_58 ();
 FILLCELL_X4 FILLER_0_12_68 ();
 FILLCELL_X1 FILLER_0_12_72 ();
 FILLCELL_X8 FILLER_0_12_90 ();
 FILLCELL_X2 FILLER_0_12_98 ();
 FILLCELL_X8 FILLER_0_12_102 ();
 FILLCELL_X1 FILLER_0_12_110 ();
 FILLCELL_X4 FILLER_0_12_114 ();
 FILLCELL_X2 FILLER_0_12_118 ();
 FILLCELL_X8 FILLER_0_12_122 ();
 FILLCELL_X2 FILLER_0_12_133 ();
 FILLCELL_X1 FILLER_0_12_135 ();
 FILLCELL_X1 FILLER_0_12_139 ();
 FILLCELL_X2 FILLER_0_12_144 ();
 FILLCELL_X1 FILLER_0_12_149 ();
 FILLCELL_X8 FILLER_0_12_153 ();
 FILLCELL_X2 FILLER_0_12_163 ();
 FILLCELL_X1 FILLER_0_12_175 ();
 FILLCELL_X1 FILLER_0_12_179 ();
 FILLCELL_X2 FILLER_0_12_187 ();
 FILLCELL_X2 FILLER_0_12_196 ();
 FILLCELL_X2 FILLER_0_12_211 ();
 FILLCELL_X1 FILLER_0_12_213 ();
 FILLCELL_X1 FILLER_0_12_216 ();
 FILLCELL_X4 FILLER_0_12_223 ();
 FILLCELL_X2 FILLER_0_12_227 ();
 FILLCELL_X1 FILLER_0_12_229 ();
 FILLCELL_X32 FILLER_0_12_233 ();
 FILLCELL_X32 FILLER_0_12_265 ();
 FILLCELL_X32 FILLER_0_12_297 ();
 FILLCELL_X32 FILLER_0_12_329 ();
 FILLCELL_X32 FILLER_0_12_361 ();
 FILLCELL_X32 FILLER_0_12_393 ();
 FILLCELL_X32 FILLER_0_12_425 ();
 FILLCELL_X8 FILLER_0_12_457 ();
 FILLCELL_X2 FILLER_0_12_465 ();
 FILLCELL_X1 FILLER_0_12_467 ();
 FILLCELL_X16 FILLER_0_13_1 ();
 FILLCELL_X8 FILLER_0_13_17 ();
 FILLCELL_X4 FILLER_0_13_25 ();
 FILLCELL_X1 FILLER_0_13_32 ();
 FILLCELL_X2 FILLER_0_13_66 ();
 FILLCELL_X8 FILLER_0_13_76 ();
 FILLCELL_X1 FILLER_0_13_84 ();
 FILLCELL_X4 FILLER_0_13_90 ();
 FILLCELL_X2 FILLER_0_13_119 ();
 FILLCELL_X4 FILLER_0_13_133 ();
 FILLCELL_X2 FILLER_0_13_141 ();
 FILLCELL_X1 FILLER_0_13_143 ();
 FILLCELL_X8 FILLER_0_13_147 ();
 FILLCELL_X4 FILLER_0_13_158 ();
 FILLCELL_X2 FILLER_0_13_162 ();
 FILLCELL_X1 FILLER_0_13_164 ();
 FILLCELL_X1 FILLER_0_13_170 ();
 FILLCELL_X2 FILLER_0_13_175 ();
 FILLCELL_X1 FILLER_0_13_177 ();
 FILLCELL_X1 FILLER_0_13_195 ();
 FILLCELL_X4 FILLER_0_13_198 ();
 FILLCELL_X8 FILLER_0_13_220 ();
 FILLCELL_X2 FILLER_0_13_228 ();
 FILLCELL_X2 FILLER_0_13_236 ();
 FILLCELL_X32 FILLER_0_13_244 ();
 FILLCELL_X32 FILLER_0_13_276 ();
 FILLCELL_X32 FILLER_0_13_308 ();
 FILLCELL_X32 FILLER_0_13_340 ();
 FILLCELL_X32 FILLER_0_13_372 ();
 FILLCELL_X32 FILLER_0_13_404 ();
 FILLCELL_X32 FILLER_0_13_436 ();
 FILLCELL_X16 FILLER_0_14_1 ();
 FILLCELL_X4 FILLER_0_14_17 ();
 FILLCELL_X2 FILLER_0_14_21 ();
 FILLCELL_X1 FILLER_0_14_23 ();
 FILLCELL_X2 FILLER_0_14_30 ();
 FILLCELL_X2 FILLER_0_14_35 ();
 FILLCELL_X1 FILLER_0_14_41 ();
 FILLCELL_X16 FILLER_0_14_45 ();
 FILLCELL_X1 FILLER_0_14_61 ();
 FILLCELL_X16 FILLER_0_14_64 ();
 FILLCELL_X4 FILLER_0_14_80 ();
 FILLCELL_X4 FILLER_0_14_91 ();
 FILLCELL_X2 FILLER_0_14_95 ();
 FILLCELL_X1 FILLER_0_14_97 ();
 FILLCELL_X2 FILLER_0_14_107 ();
 FILLCELL_X1 FILLER_0_14_109 ();
 FILLCELL_X8 FILLER_0_14_113 ();
 FILLCELL_X2 FILLER_0_14_121 ();
 FILLCELL_X1 FILLER_0_14_123 ();
 FILLCELL_X1 FILLER_0_14_127 ();
 FILLCELL_X1 FILLER_0_14_132 ();
 FILLCELL_X2 FILLER_0_14_136 ();
 FILLCELL_X2 FILLER_0_14_149 ();
 FILLCELL_X1 FILLER_0_14_155 ();
 FILLCELL_X2 FILLER_0_14_159 ();
 FILLCELL_X4 FILLER_0_14_172 ();
 FILLCELL_X2 FILLER_0_14_176 ();
 FILLCELL_X1 FILLER_0_14_178 ();
 FILLCELL_X2 FILLER_0_14_190 ();
 FILLCELL_X4 FILLER_0_14_208 ();
 FILLCELL_X1 FILLER_0_14_212 ();
 FILLCELL_X32 FILLER_0_14_235 ();
 FILLCELL_X32 FILLER_0_14_267 ();
 FILLCELL_X32 FILLER_0_14_299 ();
 FILLCELL_X32 FILLER_0_14_331 ();
 FILLCELL_X32 FILLER_0_14_363 ();
 FILLCELL_X32 FILLER_0_14_395 ();
 FILLCELL_X32 FILLER_0_14_427 ();
 FILLCELL_X8 FILLER_0_14_459 ();
 FILLCELL_X1 FILLER_0_14_467 ();
 FILLCELL_X16 FILLER_0_15_1 ();
 FILLCELL_X8 FILLER_0_15_17 ();
 FILLCELL_X1 FILLER_0_15_25 ();
 FILLCELL_X2 FILLER_0_15_33 ();
 FILLCELL_X1 FILLER_0_15_43 ();
 FILLCELL_X1 FILLER_0_15_54 ();
 FILLCELL_X1 FILLER_0_15_57 ();
 FILLCELL_X1 FILLER_0_15_61 ();
 FILLCELL_X1 FILLER_0_15_66 ();
 FILLCELL_X1 FILLER_0_15_74 ();
 FILLCELL_X8 FILLER_0_15_93 ();
 FILLCELL_X2 FILLER_0_15_101 ();
 FILLCELL_X1 FILLER_0_15_106 ();
 FILLCELL_X1 FILLER_0_15_111 ();
 FILLCELL_X1 FILLER_0_15_116 ();
 FILLCELL_X1 FILLER_0_15_121 ();
 FILLCELL_X4 FILLER_0_15_126 ();
 FILLCELL_X2 FILLER_0_15_130 ();
 FILLCELL_X1 FILLER_0_15_132 ();
 FILLCELL_X2 FILLER_0_15_137 ();
 FILLCELL_X1 FILLER_0_15_139 ();
 FILLCELL_X8 FILLER_0_15_154 ();
 FILLCELL_X4 FILLER_0_15_166 ();
 FILLCELL_X2 FILLER_0_15_170 ();
 FILLCELL_X8 FILLER_0_15_179 ();
 FILLCELL_X4 FILLER_0_15_187 ();
 FILLCELL_X2 FILLER_0_15_191 ();
 FILLCELL_X8 FILLER_0_15_225 ();
 FILLCELL_X2 FILLER_0_15_233 ();
 FILLCELL_X4 FILLER_0_15_241 ();
 FILLCELL_X2 FILLER_0_15_245 ();
 FILLCELL_X32 FILLER_0_15_249 ();
 FILLCELL_X32 FILLER_0_15_281 ();
 FILLCELL_X32 FILLER_0_15_313 ();
 FILLCELL_X32 FILLER_0_15_345 ();
 FILLCELL_X32 FILLER_0_15_377 ();
 FILLCELL_X32 FILLER_0_15_409 ();
 FILLCELL_X16 FILLER_0_15_441 ();
 FILLCELL_X8 FILLER_0_15_457 ();
 FILLCELL_X2 FILLER_0_15_465 ();
 FILLCELL_X1 FILLER_0_15_467 ();
 FILLCELL_X32 FILLER_0_16_1 ();
 FILLCELL_X4 FILLER_0_16_33 ();
 FILLCELL_X2 FILLER_0_16_49 ();
 FILLCELL_X4 FILLER_0_16_54 ();
 FILLCELL_X2 FILLER_0_16_58 ();
 FILLCELL_X1 FILLER_0_16_60 ();
 FILLCELL_X1 FILLER_0_16_64 ();
 FILLCELL_X4 FILLER_0_16_70 ();
 FILLCELL_X1 FILLER_0_16_74 ();
 FILLCELL_X8 FILLER_0_16_82 ();
 FILLCELL_X4 FILLER_0_16_90 ();
 FILLCELL_X1 FILLER_0_16_97 ();
 FILLCELL_X8 FILLER_0_16_102 ();
 FILLCELL_X2 FILLER_0_16_119 ();
 FILLCELL_X1 FILLER_0_16_121 ();
 FILLCELL_X1 FILLER_0_16_125 ();
 FILLCELL_X1 FILLER_0_16_137 ();
 FILLCELL_X2 FILLER_0_16_141 ();
 FILLCELL_X2 FILLER_0_16_147 ();
 FILLCELL_X1 FILLER_0_16_149 ();
 FILLCELL_X8 FILLER_0_16_152 ();
 FILLCELL_X1 FILLER_0_16_160 ();
 FILLCELL_X4 FILLER_0_16_167 ();
 FILLCELL_X1 FILLER_0_16_171 ();
 FILLCELL_X1 FILLER_0_16_176 ();
 FILLCELL_X2 FILLER_0_16_180 ();
 FILLCELL_X4 FILLER_0_16_188 ();
 FILLCELL_X2 FILLER_0_16_192 ();
 FILLCELL_X2 FILLER_0_16_220 ();
 FILLCELL_X8 FILLER_0_16_232 ();
 FILLCELL_X2 FILLER_0_16_240 ();
 FILLCELL_X32 FILLER_0_16_249 ();
 FILLCELL_X32 FILLER_0_16_281 ();
 FILLCELL_X32 FILLER_0_16_313 ();
 FILLCELL_X32 FILLER_0_16_345 ();
 FILLCELL_X32 FILLER_0_16_377 ();
 FILLCELL_X32 FILLER_0_16_409 ();
 FILLCELL_X16 FILLER_0_16_441 ();
 FILLCELL_X8 FILLER_0_16_457 ();
 FILLCELL_X2 FILLER_0_16_465 ();
 FILLCELL_X1 FILLER_0_16_467 ();
 FILLCELL_X16 FILLER_0_17_1 ();
 FILLCELL_X8 FILLER_0_17_17 ();
 FILLCELL_X1 FILLER_0_17_25 ();
 FILLCELL_X1 FILLER_0_17_30 ();
 FILLCELL_X1 FILLER_0_17_40 ();
 FILLCELL_X4 FILLER_0_17_52 ();
 FILLCELL_X4 FILLER_0_17_69 ();
 FILLCELL_X2 FILLER_0_17_73 ();
 FILLCELL_X1 FILLER_0_17_79 ();
 FILLCELL_X1 FILLER_0_17_83 ();
 FILLCELL_X1 FILLER_0_17_91 ();
 FILLCELL_X1 FILLER_0_17_99 ();
 FILLCELL_X2 FILLER_0_17_103 ();
 FILLCELL_X2 FILLER_0_17_108 ();
 FILLCELL_X4 FILLER_0_17_114 ();
 FILLCELL_X2 FILLER_0_17_118 ();
 FILLCELL_X1 FILLER_0_17_120 ();
 FILLCELL_X1 FILLER_0_17_124 ();
 FILLCELL_X2 FILLER_0_17_128 ();
 FILLCELL_X1 FILLER_0_17_130 ();
 FILLCELL_X2 FILLER_0_17_147 ();
 FILLCELL_X1 FILLER_0_17_149 ();
 FILLCELL_X2 FILLER_0_17_158 ();
 FILLCELL_X1 FILLER_0_17_160 ();
 FILLCELL_X4 FILLER_0_17_168 ();
 FILLCELL_X1 FILLER_0_17_172 ();
 FILLCELL_X8 FILLER_0_17_181 ();
 FILLCELL_X2 FILLER_0_17_189 ();
 FILLCELL_X8 FILLER_0_17_201 ();
 FILLCELL_X4 FILLER_0_17_209 ();
 FILLCELL_X2 FILLER_0_17_213 ();
 FILLCELL_X1 FILLER_0_17_215 ();
 FILLCELL_X4 FILLER_0_17_219 ();
 FILLCELL_X2 FILLER_0_17_223 ();
 FILLCELL_X1 FILLER_0_17_225 ();
 FILLCELL_X32 FILLER_0_17_257 ();
 FILLCELL_X32 FILLER_0_17_289 ();
 FILLCELL_X32 FILLER_0_17_321 ();
 FILLCELL_X32 FILLER_0_17_353 ();
 FILLCELL_X32 FILLER_0_17_385 ();
 FILLCELL_X32 FILLER_0_17_417 ();
 FILLCELL_X16 FILLER_0_17_449 ();
 FILLCELL_X2 FILLER_0_17_465 ();
 FILLCELL_X1 FILLER_0_17_467 ();
 FILLCELL_X16 FILLER_0_18_1 ();
 FILLCELL_X8 FILLER_0_18_17 ();
 FILLCELL_X2 FILLER_0_18_25 ();
 FILLCELL_X1 FILLER_0_18_27 ();
 FILLCELL_X1 FILLER_0_18_31 ();
 FILLCELL_X2 FILLER_0_18_37 ();
 FILLCELL_X8 FILLER_0_18_49 ();
 FILLCELL_X4 FILLER_0_18_57 ();
 FILLCELL_X4 FILLER_0_18_69 ();
 FILLCELL_X4 FILLER_0_18_88 ();
 FILLCELL_X1 FILLER_0_18_96 ();
 FILLCELL_X8 FILLER_0_18_100 ();
 FILLCELL_X4 FILLER_0_18_108 ();
 FILLCELL_X2 FILLER_0_18_112 ();
 FILLCELL_X1 FILLER_0_18_114 ();
 FILLCELL_X2 FILLER_0_18_120 ();
 FILLCELL_X1 FILLER_0_18_126 ();
 FILLCELL_X2 FILLER_0_18_131 ();
 FILLCELL_X4 FILLER_0_18_136 ();
 FILLCELL_X1 FILLER_0_18_140 ();
 FILLCELL_X4 FILLER_0_18_144 ();
 FILLCELL_X2 FILLER_0_18_151 ();
 FILLCELL_X1 FILLER_0_18_153 ();
 FILLCELL_X2 FILLER_0_18_162 ();
 FILLCELL_X1 FILLER_0_18_164 ();
 FILLCELL_X4 FILLER_0_18_172 ();
 FILLCELL_X2 FILLER_0_18_176 ();
 FILLCELL_X2 FILLER_0_18_197 ();
 FILLCELL_X1 FILLER_0_18_199 ();
 FILLCELL_X1 FILLER_0_18_210 ();
 FILLCELL_X4 FILLER_0_18_221 ();
 FILLCELL_X2 FILLER_0_18_225 ();
 FILLCELL_X4 FILLER_0_18_229 ();
 FILLCELL_X1 FILLER_0_18_233 ();
 FILLCELL_X32 FILLER_0_18_246 ();
 FILLCELL_X32 FILLER_0_18_278 ();
 FILLCELL_X32 FILLER_0_18_310 ();
 FILLCELL_X32 FILLER_0_18_342 ();
 FILLCELL_X32 FILLER_0_18_374 ();
 FILLCELL_X32 FILLER_0_18_406 ();
 FILLCELL_X16 FILLER_0_18_438 ();
 FILLCELL_X8 FILLER_0_18_454 ();
 FILLCELL_X4 FILLER_0_18_462 ();
 FILLCELL_X2 FILLER_0_18_466 ();
 FILLCELL_X8 FILLER_0_19_1 ();
 FILLCELL_X4 FILLER_0_19_9 ();
 FILLCELL_X8 FILLER_0_19_16 ();
 FILLCELL_X1 FILLER_0_19_24 ();
 FILLCELL_X4 FILLER_0_19_35 ();
 FILLCELL_X2 FILLER_0_19_39 ();
 FILLCELL_X4 FILLER_0_19_51 ();
 FILLCELL_X4 FILLER_0_19_61 ();
 FILLCELL_X1 FILLER_0_19_65 ();
 FILLCELL_X1 FILLER_0_19_74 ();
 FILLCELL_X1 FILLER_0_19_79 ();
 FILLCELL_X1 FILLER_0_19_87 ();
 FILLCELL_X2 FILLER_0_19_91 ();
 FILLCELL_X2 FILLER_0_19_97 ();
 FILLCELL_X2 FILLER_0_19_103 ();
 FILLCELL_X2 FILLER_0_19_111 ();
 FILLCELL_X8 FILLER_0_19_117 ();
 FILLCELL_X1 FILLER_0_19_132 ();
 FILLCELL_X1 FILLER_0_19_140 ();
 FILLCELL_X2 FILLER_0_19_149 ();
 FILLCELL_X4 FILLER_0_19_155 ();
 FILLCELL_X1 FILLER_0_19_162 ();
 FILLCELL_X1 FILLER_0_19_166 ();
 FILLCELL_X8 FILLER_0_19_178 ();
 FILLCELL_X16 FILLER_0_19_199 ();
 FILLCELL_X1 FILLER_0_19_215 ();
 FILLCELL_X4 FILLER_0_19_223 ();
 FILLCELL_X2 FILLER_0_19_238 ();
 FILLCELL_X32 FILLER_0_19_248 ();
 FILLCELL_X32 FILLER_0_19_280 ();
 FILLCELL_X32 FILLER_0_19_312 ();
 FILLCELL_X32 FILLER_0_19_344 ();
 FILLCELL_X32 FILLER_0_19_376 ();
 FILLCELL_X32 FILLER_0_19_408 ();
 FILLCELL_X16 FILLER_0_19_440 ();
 FILLCELL_X8 FILLER_0_19_456 ();
 FILLCELL_X4 FILLER_0_19_464 ();
 FILLCELL_X16 FILLER_0_20_1 ();
 FILLCELL_X8 FILLER_0_20_17 ();
 FILLCELL_X2 FILLER_0_20_25 ();
 FILLCELL_X1 FILLER_0_20_30 ();
 FILLCELL_X2 FILLER_0_20_34 ();
 FILLCELL_X1 FILLER_0_20_40 ();
 FILLCELL_X2 FILLER_0_20_56 ();
 FILLCELL_X1 FILLER_0_20_61 ();
 FILLCELL_X1 FILLER_0_20_65 ();
 FILLCELL_X2 FILLER_0_20_71 ();
 FILLCELL_X8 FILLER_0_20_81 ();
 FILLCELL_X2 FILLER_0_20_89 ();
 FILLCELL_X1 FILLER_0_20_91 ();
 FILLCELL_X8 FILLER_0_20_95 ();
 FILLCELL_X1 FILLER_0_20_103 ();
 FILLCELL_X2 FILLER_0_20_114 ();
 FILLCELL_X2 FILLER_0_20_125 ();
 FILLCELL_X1 FILLER_0_20_127 ();
 FILLCELL_X1 FILLER_0_20_135 ();
 FILLCELL_X2 FILLER_0_20_140 ();
 FILLCELL_X1 FILLER_0_20_142 ();
 FILLCELL_X4 FILLER_0_20_160 ();
 FILLCELL_X4 FILLER_0_20_170 ();
 FILLCELL_X1 FILLER_0_20_174 ();
 FILLCELL_X1 FILLER_0_20_179 ();
 FILLCELL_X4 FILLER_0_20_189 ();
 FILLCELL_X2 FILLER_0_20_193 ();
 FILLCELL_X16 FILLER_0_20_206 ();
 FILLCELL_X1 FILLER_0_20_222 ();
 FILLCELL_X2 FILLER_0_20_233 ();
 FILLCELL_X2 FILLER_0_20_238 ();
 FILLCELL_X1 FILLER_0_20_240 ();
 FILLCELL_X2 FILLER_0_20_244 ();
 FILLCELL_X1 FILLER_0_20_246 ();
 FILLCELL_X32 FILLER_0_20_255 ();
 FILLCELL_X32 FILLER_0_20_287 ();
 FILLCELL_X32 FILLER_0_20_319 ();
 FILLCELL_X32 FILLER_0_20_351 ();
 FILLCELL_X32 FILLER_0_20_383 ();
 FILLCELL_X32 FILLER_0_20_415 ();
 FILLCELL_X16 FILLER_0_20_447 ();
 FILLCELL_X4 FILLER_0_20_463 ();
 FILLCELL_X1 FILLER_0_20_467 ();
 FILLCELL_X16 FILLER_0_21_1 ();
 FILLCELL_X8 FILLER_0_21_17 ();
 FILLCELL_X1 FILLER_0_21_25 ();
 FILLCELL_X1 FILLER_0_21_36 ();
 FILLCELL_X2 FILLER_0_21_41 ();
 FILLCELL_X1 FILLER_0_21_49 ();
 FILLCELL_X2 FILLER_0_21_53 ();
 FILLCELL_X4 FILLER_0_21_59 ();
 FILLCELL_X2 FILLER_0_21_63 ();
 FILLCELL_X4 FILLER_0_21_71 ();
 FILLCELL_X2 FILLER_0_21_75 ();
 FILLCELL_X1 FILLER_0_21_79 ();
 FILLCELL_X4 FILLER_0_21_83 ();
 FILLCELL_X2 FILLER_0_21_97 ();
 FILLCELL_X1 FILLER_0_21_99 ();
 FILLCELL_X8 FILLER_0_21_116 ();
 FILLCELL_X4 FILLER_0_21_124 ();
 FILLCELL_X8 FILLER_0_21_142 ();
 FILLCELL_X4 FILLER_0_21_153 ();
 FILLCELL_X2 FILLER_0_21_157 ();
 FILLCELL_X1 FILLER_0_21_175 ();
 FILLCELL_X1 FILLER_0_21_201 ();
 FILLCELL_X8 FILLER_0_21_216 ();
 FILLCELL_X2 FILLER_0_21_224 ();
 FILLCELL_X32 FILLER_0_21_236 ();
 FILLCELL_X32 FILLER_0_21_268 ();
 FILLCELL_X32 FILLER_0_21_300 ();
 FILLCELL_X32 FILLER_0_21_332 ();
 FILLCELL_X32 FILLER_0_21_364 ();
 FILLCELL_X32 FILLER_0_21_396 ();
 FILLCELL_X32 FILLER_0_21_428 ();
 FILLCELL_X8 FILLER_0_21_460 ();
 FILLCELL_X16 FILLER_0_22_1 ();
 FILLCELL_X8 FILLER_0_22_17 ();
 FILLCELL_X2 FILLER_0_22_25 ();
 FILLCELL_X1 FILLER_0_22_27 ();
 FILLCELL_X8 FILLER_0_22_31 ();
 FILLCELL_X1 FILLER_0_22_39 ();
 FILLCELL_X4 FILLER_0_22_43 ();
 FILLCELL_X2 FILLER_0_22_47 ();
 FILLCELL_X1 FILLER_0_22_49 ();
 FILLCELL_X1 FILLER_0_22_53 ();
 FILLCELL_X8 FILLER_0_22_72 ();
 FILLCELL_X4 FILLER_0_22_80 ();
 FILLCELL_X2 FILLER_0_22_84 ();
 FILLCELL_X1 FILLER_0_22_86 ();
 FILLCELL_X4 FILLER_0_22_95 ();
 FILLCELL_X1 FILLER_0_22_118 ();
 FILLCELL_X1 FILLER_0_22_125 ();
 FILLCELL_X2 FILLER_0_22_133 ();
 FILLCELL_X2 FILLER_0_22_143 ();
 FILLCELL_X1 FILLER_0_22_145 ();
 FILLCELL_X2 FILLER_0_22_156 ();
 FILLCELL_X1 FILLER_0_22_158 ();
 FILLCELL_X4 FILLER_0_22_162 ();
 FILLCELL_X2 FILLER_0_22_166 ();
 FILLCELL_X1 FILLER_0_22_175 ();
 FILLCELL_X4 FILLER_0_22_179 ();
 FILLCELL_X2 FILLER_0_22_187 ();
 FILLCELL_X1 FILLER_0_22_195 ();
 FILLCELL_X2 FILLER_0_22_214 ();
 FILLCELL_X2 FILLER_0_22_229 ();
 FILLCELL_X1 FILLER_0_22_231 ();
 FILLCELL_X4 FILLER_0_22_242 ();
 FILLCELL_X32 FILLER_0_22_253 ();
 FILLCELL_X32 FILLER_0_22_285 ();
 FILLCELL_X32 FILLER_0_22_317 ();
 FILLCELL_X32 FILLER_0_22_349 ();
 FILLCELL_X32 FILLER_0_22_381 ();
 FILLCELL_X32 FILLER_0_22_413 ();
 FILLCELL_X16 FILLER_0_22_445 ();
 FILLCELL_X4 FILLER_0_22_461 ();
 FILLCELL_X2 FILLER_0_22_465 ();
 FILLCELL_X1 FILLER_0_22_467 ();
 FILLCELL_X16 FILLER_0_23_1 ();
 FILLCELL_X8 FILLER_0_23_17 ();
 FILLCELL_X1 FILLER_0_23_25 ();
 FILLCELL_X2 FILLER_0_23_29 ();
 FILLCELL_X1 FILLER_0_23_37 ();
 FILLCELL_X1 FILLER_0_23_51 ();
 FILLCELL_X1 FILLER_0_23_55 ();
 FILLCELL_X1 FILLER_0_23_63 ();
 FILLCELL_X2 FILLER_0_23_68 ();
 FILLCELL_X2 FILLER_0_23_94 ();
 FILLCELL_X2 FILLER_0_23_100 ();
 FILLCELL_X1 FILLER_0_23_102 ();
 FILLCELL_X4 FILLER_0_23_112 ();
 FILLCELL_X1 FILLER_0_23_116 ();
 FILLCELL_X4 FILLER_0_23_129 ();
 FILLCELL_X1 FILLER_0_23_133 ();
 FILLCELL_X4 FILLER_0_23_138 ();
 FILLCELL_X1 FILLER_0_23_142 ();
 FILLCELL_X2 FILLER_0_23_153 ();
 FILLCELL_X1 FILLER_0_23_155 ();
 FILLCELL_X1 FILLER_0_23_159 ();
 FILLCELL_X4 FILLER_0_23_234 ();
 FILLCELL_X2 FILLER_0_23_238 ();
 FILLCELL_X4 FILLER_0_23_243 ();
 FILLCELL_X2 FILLER_0_23_247 ();
 FILLCELL_X1 FILLER_0_23_255 ();
 FILLCELL_X32 FILLER_0_23_260 ();
 FILLCELL_X32 FILLER_0_23_292 ();
 FILLCELL_X32 FILLER_0_23_324 ();
 FILLCELL_X32 FILLER_0_23_356 ();
 FILLCELL_X32 FILLER_0_23_388 ();
 FILLCELL_X32 FILLER_0_23_420 ();
 FILLCELL_X16 FILLER_0_23_452 ();
 FILLCELL_X8 FILLER_0_24_1 ();
 FILLCELL_X16 FILLER_0_24_12 ();
 FILLCELL_X2 FILLER_0_24_31 ();
 FILLCELL_X2 FILLER_0_24_36 ();
 FILLCELL_X2 FILLER_0_24_41 ();
 FILLCELL_X4 FILLER_0_24_54 ();
 FILLCELL_X1 FILLER_0_24_58 ();
 FILLCELL_X8 FILLER_0_24_62 ();
 FILLCELL_X4 FILLER_0_24_70 ();
 FILLCELL_X1 FILLER_0_24_74 ();
 FILLCELL_X4 FILLER_0_24_78 ();
 FILLCELL_X2 FILLER_0_24_82 ();
 FILLCELL_X1 FILLER_0_24_84 ();
 FILLCELL_X1 FILLER_0_24_98 ();
 FILLCELL_X2 FILLER_0_24_107 ();
 FILLCELL_X2 FILLER_0_24_113 ();
 FILLCELL_X8 FILLER_0_24_135 ();
 FILLCELL_X2 FILLER_0_24_143 ();
 FILLCELL_X1 FILLER_0_24_145 ();
 FILLCELL_X2 FILLER_0_24_150 ();
 FILLCELL_X1 FILLER_0_24_152 ();
 FILLCELL_X1 FILLER_0_24_155 ();
 FILLCELL_X8 FILLER_0_24_159 ();
 FILLCELL_X2 FILLER_0_24_187 ();
 FILLCELL_X1 FILLER_0_24_189 ();
 FILLCELL_X1 FILLER_0_24_193 ();
 FILLCELL_X16 FILLER_0_24_197 ();
 FILLCELL_X8 FILLER_0_24_213 ();
 FILLCELL_X4 FILLER_0_24_221 ();
 FILLCELL_X1 FILLER_0_24_247 ();
 FILLCELL_X32 FILLER_0_24_254 ();
 FILLCELL_X32 FILLER_0_24_286 ();
 FILLCELL_X32 FILLER_0_24_318 ();
 FILLCELL_X32 FILLER_0_24_350 ();
 FILLCELL_X32 FILLER_0_24_382 ();
 FILLCELL_X32 FILLER_0_24_414 ();
 FILLCELL_X16 FILLER_0_24_446 ();
 FILLCELL_X4 FILLER_0_24_462 ();
 FILLCELL_X2 FILLER_0_24_466 ();
 FILLCELL_X8 FILLER_0_25_1 ();
 FILLCELL_X4 FILLER_0_25_9 ();
 FILLCELL_X2 FILLER_0_25_13 ();
 FILLCELL_X1 FILLER_0_25_15 ();
 FILLCELL_X16 FILLER_0_25_18 ();
 FILLCELL_X8 FILLER_0_25_34 ();
 FILLCELL_X2 FILLER_0_25_42 ();
 FILLCELL_X1 FILLER_0_25_44 ();
 FILLCELL_X1 FILLER_0_25_54 ();
 FILLCELL_X4 FILLER_0_25_69 ();
 FILLCELL_X2 FILLER_0_25_73 ();
 FILLCELL_X1 FILLER_0_25_75 ();
 FILLCELL_X4 FILLER_0_25_80 ();
 FILLCELL_X1 FILLER_0_25_84 ();
 FILLCELL_X2 FILLER_0_25_111 ();
 FILLCELL_X1 FILLER_0_25_113 ();
 FILLCELL_X4 FILLER_0_25_117 ();
 FILLCELL_X2 FILLER_0_25_129 ();
 FILLCELL_X8 FILLER_0_25_141 ();
 FILLCELL_X4 FILLER_0_25_149 ();
 FILLCELL_X4 FILLER_0_25_161 ();
 FILLCELL_X1 FILLER_0_25_174 ();
 FILLCELL_X1 FILLER_0_25_178 ();
 FILLCELL_X8 FILLER_0_25_205 ();
 FILLCELL_X4 FILLER_0_25_213 ();
 FILLCELL_X2 FILLER_0_25_217 ();
 FILLCELL_X1 FILLER_0_25_219 ();
 FILLCELL_X2 FILLER_0_25_222 ();
 FILLCELL_X1 FILLER_0_25_224 ();
 FILLCELL_X2 FILLER_0_25_235 ();
 FILLCELL_X1 FILLER_0_25_239 ();
 FILLCELL_X1 FILLER_0_25_247 ();
 FILLCELL_X2 FILLER_0_25_269 ();
 FILLCELL_X1 FILLER_0_25_271 ();
 FILLCELL_X1 FILLER_0_25_275 ();
 FILLCELL_X1 FILLER_0_25_282 ();
 FILLCELL_X2 FILLER_0_25_286 ();
 FILLCELL_X8 FILLER_0_25_291 ();
 FILLCELL_X2 FILLER_0_25_299 ();
 FILLCELL_X1 FILLER_0_25_304 ();
 FILLCELL_X2 FILLER_0_25_308 ();
 FILLCELL_X4 FILLER_0_25_312 ();
 FILLCELL_X2 FILLER_0_25_319 ();
 FILLCELL_X1 FILLER_0_25_324 ();
 FILLCELL_X2 FILLER_0_25_336 ();
 FILLCELL_X2 FILLER_0_25_343 ();
 FILLCELL_X1 FILLER_0_25_345 ();
 FILLCELL_X16 FILLER_0_25_352 ();
 FILLCELL_X1 FILLER_0_25_368 ();
 FILLCELL_X1 FILLER_0_25_378 ();
 FILLCELL_X8 FILLER_0_25_381 ();
 FILLCELL_X2 FILLER_0_25_389 ();
 FILLCELL_X1 FILLER_0_25_391 ();
 FILLCELL_X32 FILLER_0_25_397 ();
 FILLCELL_X32 FILLER_0_25_429 ();
 FILLCELL_X4 FILLER_0_25_461 ();
 FILLCELL_X2 FILLER_0_25_465 ();
 FILLCELL_X1 FILLER_0_25_467 ();
 FILLCELL_X32 FILLER_0_26_1 ();
 FILLCELL_X2 FILLER_0_26_33 ();
 FILLCELL_X4 FILLER_0_26_49 ();
 FILLCELL_X1 FILLER_0_26_53 ();
 FILLCELL_X16 FILLER_0_26_56 ();
 FILLCELL_X2 FILLER_0_26_72 ();
 FILLCELL_X1 FILLER_0_26_74 ();
 FILLCELL_X2 FILLER_0_26_80 ();
 FILLCELL_X1 FILLER_0_26_82 ();
 FILLCELL_X2 FILLER_0_26_86 ();
 FILLCELL_X1 FILLER_0_26_88 ();
 FILLCELL_X2 FILLER_0_26_92 ();
 FILLCELL_X1 FILLER_0_26_97 ();
 FILLCELL_X4 FILLER_0_26_102 ();
 FILLCELL_X2 FILLER_0_26_106 ();
 FILLCELL_X1 FILLER_0_26_108 ();
 FILLCELL_X1 FILLER_0_26_116 ();
 FILLCELL_X4 FILLER_0_26_125 ();
 FILLCELL_X1 FILLER_0_26_129 ();
 FILLCELL_X2 FILLER_0_26_133 ();
 FILLCELL_X1 FILLER_0_26_138 ();
 FILLCELL_X2 FILLER_0_26_149 ();
 FILLCELL_X1 FILLER_0_26_151 ();
 FILLCELL_X1 FILLER_0_26_155 ();
 FILLCELL_X2 FILLER_0_26_160 ();
 FILLCELL_X1 FILLER_0_26_162 ();
 FILLCELL_X2 FILLER_0_26_169 ();
 FILLCELL_X8 FILLER_0_26_179 ();
 FILLCELL_X2 FILLER_0_26_187 ();
 FILLCELL_X1 FILLER_0_26_189 ();
 FILLCELL_X2 FILLER_0_26_200 ();
 FILLCELL_X1 FILLER_0_26_217 ();
 FILLCELL_X2 FILLER_0_26_224 ();
 FILLCELL_X2 FILLER_0_26_236 ();
 FILLCELL_X1 FILLER_0_26_238 ();
 FILLCELL_X2 FILLER_0_26_249 ();
 FILLCELL_X1 FILLER_0_26_251 ();
 FILLCELL_X4 FILLER_0_26_262 ();
 FILLCELL_X2 FILLER_0_26_266 ();
 FILLCELL_X2 FILLER_0_26_282 ();
 FILLCELL_X2 FILLER_0_26_293 ();
 FILLCELL_X1 FILLER_0_26_295 ();
 FILLCELL_X4 FILLER_0_26_304 ();
 FILLCELL_X2 FILLER_0_26_318 ();
 FILLCELL_X2 FILLER_0_26_327 ();
 FILLCELL_X4 FILLER_0_26_333 ();
 FILLCELL_X1 FILLER_0_26_337 ();
 FILLCELL_X2 FILLER_0_26_372 ();
 FILLCELL_X1 FILLER_0_26_385 ();
 FILLCELL_X2 FILLER_0_26_389 ();
 FILLCELL_X1 FILLER_0_26_395 ();
 FILLCELL_X2 FILLER_0_26_399 ();
 FILLCELL_X2 FILLER_0_26_407 ();
 FILLCELL_X1 FILLER_0_26_414 ();
 FILLCELL_X16 FILLER_0_26_448 ();
 FILLCELL_X4 FILLER_0_26_464 ();
 FILLCELL_X16 FILLER_0_27_1 ();
 FILLCELL_X16 FILLER_0_27_20 ();
 FILLCELL_X4 FILLER_0_27_36 ();
 FILLCELL_X1 FILLER_0_27_43 ();
 FILLCELL_X1 FILLER_0_27_57 ();
 FILLCELL_X1 FILLER_0_27_64 ();
 FILLCELL_X4 FILLER_0_27_69 ();
 FILLCELL_X2 FILLER_0_27_78 ();
 FILLCELL_X1 FILLER_0_27_87 ();
 FILLCELL_X1 FILLER_0_27_92 ();
 FILLCELL_X8 FILLER_0_27_95 ();
 FILLCELL_X4 FILLER_0_27_111 ();
 FILLCELL_X2 FILLER_0_27_117 ();
 FILLCELL_X2 FILLER_0_27_126 ();
 FILLCELL_X4 FILLER_0_27_133 ();
 FILLCELL_X1 FILLER_0_27_156 ();
 FILLCELL_X8 FILLER_0_27_159 ();
 FILLCELL_X2 FILLER_0_27_167 ();
 FILLCELL_X1 FILLER_0_27_169 ();
 FILLCELL_X4 FILLER_0_27_174 ();
 FILLCELL_X1 FILLER_0_27_178 ();
 FILLCELL_X4 FILLER_0_27_183 ();
 FILLCELL_X8 FILLER_0_27_197 ();
 FILLCELL_X4 FILLER_0_27_205 ();
 FILLCELL_X2 FILLER_0_27_209 ();
 FILLCELL_X1 FILLER_0_27_211 ();
 FILLCELL_X2 FILLER_0_27_216 ();
 FILLCELL_X8 FILLER_0_27_231 ();
 FILLCELL_X2 FILLER_0_27_239 ();
 FILLCELL_X16 FILLER_0_27_247 ();
 FILLCELL_X4 FILLER_0_27_263 ();
 FILLCELL_X8 FILLER_0_27_270 ();
 FILLCELL_X2 FILLER_0_27_278 ();
 FILLCELL_X1 FILLER_0_27_280 ();
 FILLCELL_X8 FILLER_0_27_284 ();
 FILLCELL_X2 FILLER_0_27_292 ();
 FILLCELL_X1 FILLER_0_27_294 ();
 FILLCELL_X2 FILLER_0_27_306 ();
 FILLCELL_X2 FILLER_0_27_315 ();
 FILLCELL_X1 FILLER_0_27_317 ();
 FILLCELL_X1 FILLER_0_27_322 ();
 FILLCELL_X4 FILLER_0_27_327 ();
 FILLCELL_X1 FILLER_0_27_331 ();
 FILLCELL_X8 FILLER_0_27_339 ();
 FILLCELL_X4 FILLER_0_27_347 ();
 FILLCELL_X8 FILLER_0_27_365 ();
 FILLCELL_X4 FILLER_0_27_373 ();
 FILLCELL_X2 FILLER_0_27_381 ();
 FILLCELL_X2 FILLER_0_27_387 ();
 FILLCELL_X1 FILLER_0_27_389 ();
 FILLCELL_X2 FILLER_0_27_393 ();
 FILLCELL_X1 FILLER_0_27_395 ();
 FILLCELL_X1 FILLER_0_27_400 ();
 FILLCELL_X2 FILLER_0_27_405 ();
 FILLCELL_X1 FILLER_0_27_410 ();
 FILLCELL_X2 FILLER_0_27_415 ();
 FILLCELL_X2 FILLER_0_27_420 ();
 FILLCELL_X4 FILLER_0_27_427 ();
 FILLCELL_X1 FILLER_0_27_431 ();
 FILLCELL_X16 FILLER_0_27_449 ();
 FILLCELL_X2 FILLER_0_27_465 ();
 FILLCELL_X1 FILLER_0_27_467 ();
 FILLCELL_X32 FILLER_0_28_4 ();
 FILLCELL_X8 FILLER_0_28_36 ();
 FILLCELL_X1 FILLER_0_28_44 ();
 FILLCELL_X2 FILLER_0_28_48 ();
 FILLCELL_X1 FILLER_0_28_55 ();
 FILLCELL_X2 FILLER_0_28_61 ();
 FILLCELL_X4 FILLER_0_28_65 ();
 FILLCELL_X2 FILLER_0_28_69 ();
 FILLCELL_X2 FILLER_0_28_73 ();
 FILLCELL_X1 FILLER_0_28_75 ();
 FILLCELL_X2 FILLER_0_28_83 ();
 FILLCELL_X1 FILLER_0_28_119 ();
 FILLCELL_X2 FILLER_0_28_124 ();
 FILLCELL_X1 FILLER_0_28_126 ();
 FILLCELL_X4 FILLER_0_28_139 ();
 FILLCELL_X2 FILLER_0_28_143 ();
 FILLCELL_X1 FILLER_0_28_157 ();
 FILLCELL_X8 FILLER_0_28_173 ();
 FILLCELL_X4 FILLER_0_28_187 ();
 FILLCELL_X2 FILLER_0_28_191 ();
 FILLCELL_X2 FILLER_0_28_202 ();
 FILLCELL_X1 FILLER_0_28_204 ();
 FILLCELL_X1 FILLER_0_28_228 ();
 FILLCELL_X8 FILLER_0_28_235 ();
 FILLCELL_X4 FILLER_0_28_243 ();
 FILLCELL_X2 FILLER_0_28_247 ();
 FILLCELL_X8 FILLER_0_28_252 ();
 FILLCELL_X1 FILLER_0_28_260 ();
 FILLCELL_X1 FILLER_0_28_275 ();
 FILLCELL_X2 FILLER_0_28_287 ();
 FILLCELL_X1 FILLER_0_28_298 ();
 FILLCELL_X1 FILLER_0_28_301 ();
 FILLCELL_X1 FILLER_0_28_310 ();
 FILLCELL_X2 FILLER_0_28_314 ();
 FILLCELL_X8 FILLER_0_28_323 ();
 FILLCELL_X1 FILLER_0_28_331 ();
 FILLCELL_X4 FILLER_0_28_339 ();
 FILLCELL_X2 FILLER_0_28_343 ();
 FILLCELL_X4 FILLER_0_28_348 ();
 FILLCELL_X4 FILLER_0_28_358 ();
 FILLCELL_X1 FILLER_0_28_362 ();
 FILLCELL_X1 FILLER_0_28_367 ();
 FILLCELL_X1 FILLER_0_28_372 ();
 FILLCELL_X2 FILLER_0_28_377 ();
 FILLCELL_X1 FILLER_0_28_379 ();
 FILLCELL_X2 FILLER_0_28_383 ();
 FILLCELL_X4 FILLER_0_28_393 ();
 FILLCELL_X2 FILLER_0_28_409 ();
 FILLCELL_X2 FILLER_0_28_414 ();
 FILLCELL_X1 FILLER_0_28_416 ();
 FILLCELL_X1 FILLER_0_28_424 ();
 FILLCELL_X4 FILLER_0_28_428 ();
 FILLCELL_X2 FILLER_0_28_432 ();
 FILLCELL_X1 FILLER_0_28_434 ();
 FILLCELL_X2 FILLER_0_28_438 ();
 FILLCELL_X16 FILLER_0_28_446 ();
 FILLCELL_X4 FILLER_0_28_462 ();
 FILLCELL_X2 FILLER_0_28_466 ();
 FILLCELL_X4 FILLER_0_29_4 ();
 FILLCELL_X1 FILLER_0_29_8 ();
 FILLCELL_X4 FILLER_0_29_15 ();
 FILLCELL_X4 FILLER_0_29_22 ();
 FILLCELL_X1 FILLER_0_29_26 ();
 FILLCELL_X8 FILLER_0_29_30 ();
 FILLCELL_X4 FILLER_0_29_38 ();
 FILLCELL_X2 FILLER_0_29_42 ();
 FILLCELL_X16 FILLER_0_29_48 ();
 FILLCELL_X2 FILLER_0_29_64 ();
 FILLCELL_X1 FILLER_0_29_66 ();
 FILLCELL_X8 FILLER_0_29_69 ();
 FILLCELL_X4 FILLER_0_29_77 ();
 FILLCELL_X2 FILLER_0_29_85 ();
 FILLCELL_X4 FILLER_0_29_94 ();
 FILLCELL_X1 FILLER_0_29_98 ();
 FILLCELL_X4 FILLER_0_29_108 ();
 FILLCELL_X1 FILLER_0_29_112 ();
 FILLCELL_X16 FILLER_0_29_117 ();
 FILLCELL_X2 FILLER_0_29_166 ();
 FILLCELL_X4 FILLER_0_29_178 ();
 FILLCELL_X8 FILLER_0_29_211 ();
 FILLCELL_X1 FILLER_0_29_219 ();
 FILLCELL_X8 FILLER_0_29_223 ();
 FILLCELL_X8 FILLER_0_29_236 ();
 FILLCELL_X4 FILLER_0_29_244 ();
 FILLCELL_X2 FILLER_0_29_248 ();
 FILLCELL_X4 FILLER_0_29_260 ();
 FILLCELL_X1 FILLER_0_29_264 ();
 FILLCELL_X1 FILLER_0_29_276 ();
 FILLCELL_X8 FILLER_0_29_289 ();
 FILLCELL_X4 FILLER_0_29_297 ();
 FILLCELL_X2 FILLER_0_29_301 ();
 FILLCELL_X1 FILLER_0_29_303 ();
 FILLCELL_X4 FILLER_0_29_311 ();
 FILLCELL_X1 FILLER_0_29_315 ();
 FILLCELL_X4 FILLER_0_29_330 ();
 FILLCELL_X1 FILLER_0_29_334 ();
 FILLCELL_X2 FILLER_0_29_343 ();
 FILLCELL_X4 FILLER_0_29_355 ();
 FILLCELL_X2 FILLER_0_29_359 ();
 FILLCELL_X2 FILLER_0_29_364 ();
 FILLCELL_X4 FILLER_0_29_370 ();
 FILLCELL_X1 FILLER_0_29_376 ();
 FILLCELL_X4 FILLER_0_29_380 ();
 FILLCELL_X1 FILLER_0_29_384 ();
 FILLCELL_X4 FILLER_0_29_391 ();
 FILLCELL_X1 FILLER_0_29_395 ();
 FILLCELL_X4 FILLER_0_29_402 ();
 FILLCELL_X1 FILLER_0_29_406 ();
 FILLCELL_X2 FILLER_0_29_421 ();
 FILLCELL_X4 FILLER_0_29_427 ();
 FILLCELL_X2 FILLER_0_29_431 ();
 FILLCELL_X1 FILLER_0_29_433 ();
 FILLCELL_X1 FILLER_0_29_438 ();
 FILLCELL_X16 FILLER_0_29_447 ();
 FILLCELL_X4 FILLER_0_29_463 ();
 FILLCELL_X1 FILLER_0_29_467 ();
 FILLCELL_X2 FILLER_0_30_17 ();
 FILLCELL_X1 FILLER_0_30_22 ();
 FILLCELL_X1 FILLER_0_30_32 ();
 FILLCELL_X2 FILLER_0_30_42 ();
 FILLCELL_X2 FILLER_0_30_54 ();
 FILLCELL_X1 FILLER_0_30_56 ();
 FILLCELL_X2 FILLER_0_30_64 ();
 FILLCELL_X2 FILLER_0_30_73 ();
 FILLCELL_X1 FILLER_0_30_75 ();
 FILLCELL_X8 FILLER_0_30_108 ();
 FILLCELL_X8 FILLER_0_30_124 ();
 FILLCELL_X2 FILLER_0_30_132 ();
 FILLCELL_X1 FILLER_0_30_138 ();
 FILLCELL_X1 FILLER_0_30_149 ();
 FILLCELL_X2 FILLER_0_30_172 ();
 FILLCELL_X4 FILLER_0_30_224 ();
 FILLCELL_X1 FILLER_0_30_228 ();
 FILLCELL_X2 FILLER_0_30_236 ();
 FILLCELL_X1 FILLER_0_30_257 ();
 FILLCELL_X1 FILLER_0_30_261 ();
 FILLCELL_X16 FILLER_0_30_269 ();
 FILLCELL_X2 FILLER_0_30_285 ();
 FILLCELL_X1 FILLER_0_30_287 ();
 FILLCELL_X1 FILLER_0_30_298 ();
 FILLCELL_X4 FILLER_0_30_310 ();
 FILLCELL_X2 FILLER_0_30_314 ();
 FILLCELL_X1 FILLER_0_30_316 ();
 FILLCELL_X8 FILLER_0_30_321 ();
 FILLCELL_X2 FILLER_0_30_329 ();
 FILLCELL_X1 FILLER_0_30_331 ();
 FILLCELL_X2 FILLER_0_30_339 ();
 FILLCELL_X1 FILLER_0_30_341 ();
 FILLCELL_X4 FILLER_0_30_350 ();
 FILLCELL_X1 FILLER_0_30_354 ();
 FILLCELL_X2 FILLER_0_30_359 ();
 FILLCELL_X1 FILLER_0_30_361 ();
 FILLCELL_X1 FILLER_0_30_366 ();
 FILLCELL_X4 FILLER_0_30_380 ();
 FILLCELL_X2 FILLER_0_30_384 ();
 FILLCELL_X1 FILLER_0_30_386 ();
 FILLCELL_X1 FILLER_0_30_397 ();
 FILLCELL_X1 FILLER_0_30_402 ();
 FILLCELL_X1 FILLER_0_30_423 ();
 FILLCELL_X2 FILLER_0_30_436 ();
 FILLCELL_X16 FILLER_0_30_442 ();
 FILLCELL_X8 FILLER_0_30_458 ();
 FILLCELL_X2 FILLER_0_30_466 ();
 FILLCELL_X1 FILLER_0_31_1 ();
 FILLCELL_X2 FILLER_0_31_38 ();
 FILLCELL_X1 FILLER_0_31_40 ();
 FILLCELL_X2 FILLER_0_31_47 ();
 FILLCELL_X8 FILLER_0_31_59 ();
 FILLCELL_X2 FILLER_0_31_67 ();
 FILLCELL_X1 FILLER_0_31_79 ();
 FILLCELL_X1 FILLER_0_31_85 ();
 FILLCELL_X1 FILLER_0_31_89 ();
 FILLCELL_X2 FILLER_0_31_93 ();
 FILLCELL_X1 FILLER_0_31_95 ();
 FILLCELL_X4 FILLER_0_31_99 ();
 FILLCELL_X1 FILLER_0_31_103 ();
 FILLCELL_X4 FILLER_0_31_117 ();
 FILLCELL_X1 FILLER_0_31_121 ();
 FILLCELL_X4 FILLER_0_31_132 ();
 FILLCELL_X2 FILLER_0_31_136 ();
 FILLCELL_X4 FILLER_0_31_145 ();
 FILLCELL_X2 FILLER_0_31_149 ();
 FILLCELL_X1 FILLER_0_31_155 ();
 FILLCELL_X4 FILLER_0_31_159 ();
 FILLCELL_X2 FILLER_0_31_163 ();
 FILLCELL_X1 FILLER_0_31_165 ();
 FILLCELL_X2 FILLER_0_31_175 ();
 FILLCELL_X8 FILLER_0_31_183 ();
 FILLCELL_X2 FILLER_0_31_202 ();
 FILLCELL_X8 FILLER_0_31_214 ();
 FILLCELL_X4 FILLER_0_31_222 ();
 FILLCELL_X2 FILLER_0_31_226 ();
 FILLCELL_X4 FILLER_0_31_238 ();
 FILLCELL_X2 FILLER_0_31_242 ();
 FILLCELL_X4 FILLER_0_31_250 ();
 FILLCELL_X2 FILLER_0_31_254 ();
 FILLCELL_X2 FILLER_0_31_260 ();
 FILLCELL_X2 FILLER_0_31_269 ();
 FILLCELL_X4 FILLER_0_31_284 ();
 FILLCELL_X2 FILLER_0_31_288 ();
 FILLCELL_X4 FILLER_0_31_294 ();
 FILLCELL_X1 FILLER_0_31_301 ();
 FILLCELL_X8 FILLER_0_31_309 ();
 FILLCELL_X2 FILLER_0_31_320 ();
 FILLCELL_X1 FILLER_0_31_322 ();
 FILLCELL_X2 FILLER_0_31_346 ();
 FILLCELL_X1 FILLER_0_31_348 ();
 FILLCELL_X1 FILLER_0_31_352 ();
 FILLCELL_X2 FILLER_0_31_360 ();
 FILLCELL_X2 FILLER_0_31_373 ();
 FILLCELL_X1 FILLER_0_31_400 ();
 FILLCELL_X2 FILLER_0_31_404 ();
 FILLCELL_X1 FILLER_0_31_409 ();
 FILLCELL_X4 FILLER_0_31_418 ();
 FILLCELL_X2 FILLER_0_31_425 ();
 FILLCELL_X2 FILLER_0_31_430 ();
 FILLCELL_X2 FILLER_0_31_436 ();
 FILLCELL_X16 FILLER_0_31_450 ();
 FILLCELL_X2 FILLER_0_31_466 ();
 FILLCELL_X2 FILLER_0_32_1 ();
 FILLCELL_X1 FILLER_0_32_3 ();
 FILLCELL_X1 FILLER_0_32_11 ();
 FILLCELL_X1 FILLER_0_32_14 ();
 FILLCELL_X2 FILLER_0_32_18 ();
 FILLCELL_X8 FILLER_0_32_23 ();
 FILLCELL_X4 FILLER_0_32_41 ();
 FILLCELL_X1 FILLER_0_32_45 ();
 FILLCELL_X1 FILLER_0_32_50 ();
 FILLCELL_X1 FILLER_0_32_57 ();
 FILLCELL_X4 FILLER_0_32_65 ();
 FILLCELL_X2 FILLER_0_32_74 ();
 FILLCELL_X1 FILLER_0_32_76 ();
 FILLCELL_X4 FILLER_0_32_81 ();
 FILLCELL_X2 FILLER_0_32_85 ();
 FILLCELL_X1 FILLER_0_32_87 ();
 FILLCELL_X1 FILLER_0_32_97 ();
 FILLCELL_X1 FILLER_0_32_102 ();
 FILLCELL_X1 FILLER_0_32_106 ();
 FILLCELL_X1 FILLER_0_32_110 ();
 FILLCELL_X2 FILLER_0_32_116 ();
 FILLCELL_X2 FILLER_0_32_130 ();
 FILLCELL_X1 FILLER_0_32_132 ();
 FILLCELL_X4 FILLER_0_32_145 ();
 FILLCELL_X2 FILLER_0_32_149 ();
 FILLCELL_X1 FILLER_0_32_164 ();
 FILLCELL_X1 FILLER_0_32_168 ();
 FILLCELL_X1 FILLER_0_32_172 ();
 FILLCELL_X2 FILLER_0_32_179 ();
 FILLCELL_X2 FILLER_0_32_195 ();
 FILLCELL_X2 FILLER_0_32_215 ();
 FILLCELL_X1 FILLER_0_32_217 ();
 FILLCELL_X1 FILLER_0_32_224 ();
 FILLCELL_X2 FILLER_0_32_233 ();
 FILLCELL_X1 FILLER_0_32_235 ();
 FILLCELL_X2 FILLER_0_32_239 ();
 FILLCELL_X2 FILLER_0_32_256 ();
 FILLCELL_X1 FILLER_0_32_258 ();
 FILLCELL_X1 FILLER_0_32_262 ();
 FILLCELL_X2 FILLER_0_32_283 ();
 FILLCELL_X1 FILLER_0_32_292 ();
 FILLCELL_X4 FILLER_0_32_300 ();
 FILLCELL_X1 FILLER_0_32_304 ();
 FILLCELL_X2 FILLER_0_32_309 ();
 FILLCELL_X1 FILLER_0_32_311 ();
 FILLCELL_X8 FILLER_0_32_317 ();
 FILLCELL_X1 FILLER_0_32_325 ();
 FILLCELL_X4 FILLER_0_32_329 ();
 FILLCELL_X4 FILLER_0_32_335 ();
 FILLCELL_X2 FILLER_0_32_339 ();
 FILLCELL_X1 FILLER_0_32_341 ();
 FILLCELL_X4 FILLER_0_32_346 ();
 FILLCELL_X1 FILLER_0_32_350 ();
 FILLCELL_X8 FILLER_0_32_355 ();
 FILLCELL_X4 FILLER_0_32_363 ();
 FILLCELL_X2 FILLER_0_32_367 ();
 FILLCELL_X8 FILLER_0_32_372 ();
 FILLCELL_X2 FILLER_0_32_380 ();
 FILLCELL_X2 FILLER_0_32_386 ();
 FILLCELL_X1 FILLER_0_32_388 ();
 FILLCELL_X1 FILLER_0_32_391 ();
 FILLCELL_X2 FILLER_0_32_418 ();
 FILLCELL_X4 FILLER_0_32_422 ();
 FILLCELL_X4 FILLER_0_32_433 ();
 FILLCELL_X2 FILLER_0_32_440 ();
 FILLCELL_X16 FILLER_0_32_452 ();
 FILLCELL_X2 FILLER_0_33_16 ();
 FILLCELL_X8 FILLER_0_33_21 ();
 FILLCELL_X1 FILLER_0_33_29 ();
 FILLCELL_X4 FILLER_0_33_33 ();
 FILLCELL_X2 FILLER_0_33_40 ();
 FILLCELL_X2 FILLER_0_33_55 ();
 FILLCELL_X2 FILLER_0_33_62 ();
 FILLCELL_X1 FILLER_0_33_64 ();
 FILLCELL_X2 FILLER_0_33_72 ();
 FILLCELL_X4 FILLER_0_33_105 ();
 FILLCELL_X1 FILLER_0_33_109 ();
 FILLCELL_X1 FILLER_0_33_117 ();
 FILLCELL_X1 FILLER_0_33_128 ();
 FILLCELL_X1 FILLER_0_33_138 ();
 FILLCELL_X1 FILLER_0_33_145 ();
 FILLCELL_X2 FILLER_0_33_156 ();
 FILLCELL_X1 FILLER_0_33_201 ();
 FILLCELL_X16 FILLER_0_33_206 ();
 FILLCELL_X2 FILLER_0_33_222 ();
 FILLCELL_X1 FILLER_0_33_224 ();
 FILLCELL_X4 FILLER_0_33_232 ();
 FILLCELL_X2 FILLER_0_33_236 ();
 FILLCELL_X1 FILLER_0_33_238 ();
 FILLCELL_X2 FILLER_0_33_243 ();
 FILLCELL_X1 FILLER_0_33_245 ();
 FILLCELL_X1 FILLER_0_33_249 ();
 FILLCELL_X2 FILLER_0_33_255 ();
 FILLCELL_X2 FILLER_0_33_262 ();
 FILLCELL_X2 FILLER_0_33_271 ();
 FILLCELL_X1 FILLER_0_33_286 ();
 FILLCELL_X2 FILLER_0_33_292 ();
 FILLCELL_X1 FILLER_0_33_294 ();
 FILLCELL_X16 FILLER_0_33_298 ();
 FILLCELL_X2 FILLER_0_33_314 ();
 FILLCELL_X1 FILLER_0_33_320 ();
 FILLCELL_X8 FILLER_0_33_327 ();
 FILLCELL_X1 FILLER_0_33_335 ();
 FILLCELL_X8 FILLER_0_33_347 ();
 FILLCELL_X1 FILLER_0_33_367 ();
 FILLCELL_X2 FILLER_0_33_379 ();
 FILLCELL_X4 FILLER_0_33_391 ();
 FILLCELL_X2 FILLER_0_33_398 ();
 FILLCELL_X1 FILLER_0_33_407 ();
 FILLCELL_X1 FILLER_0_33_411 ();
 FILLCELL_X2 FILLER_0_33_420 ();
 FILLCELL_X2 FILLER_0_33_430 ();
 FILLCELL_X1 FILLER_0_33_432 ();
 FILLCELL_X4 FILLER_0_33_436 ();
 FILLCELL_X2 FILLER_0_33_440 ();
 FILLCELL_X1 FILLER_0_33_442 ();
 FILLCELL_X8 FILLER_0_33_453 ();
 FILLCELL_X4 FILLER_0_33_461 ();
 FILLCELL_X2 FILLER_0_33_465 ();
 FILLCELL_X1 FILLER_0_33_467 ();
 FILLCELL_X4 FILLER_0_34_1 ();
 FILLCELL_X8 FILLER_0_34_8 ();
 FILLCELL_X2 FILLER_0_34_16 ();
 FILLCELL_X4 FILLER_0_34_21 ();
 FILLCELL_X2 FILLER_0_34_25 ();
 FILLCELL_X2 FILLER_0_34_34 ();
 FILLCELL_X1 FILLER_0_34_42 ();
 FILLCELL_X4 FILLER_0_34_51 ();
 FILLCELL_X1 FILLER_0_34_55 ();
 FILLCELL_X8 FILLER_0_34_59 ();
 FILLCELL_X2 FILLER_0_34_67 ();
 FILLCELL_X1 FILLER_0_34_73 ();
 FILLCELL_X1 FILLER_0_34_77 ();
 FILLCELL_X4 FILLER_0_34_85 ();
 FILLCELL_X2 FILLER_0_34_89 ();
 FILLCELL_X1 FILLER_0_34_91 ();
 FILLCELL_X4 FILLER_0_34_94 ();
 FILLCELL_X8 FILLER_0_34_100 ();
 FILLCELL_X2 FILLER_0_34_108 ();
 FILLCELL_X1 FILLER_0_34_110 ();
 FILLCELL_X4 FILLER_0_34_118 ();
 FILLCELL_X2 FILLER_0_34_132 ();
 FILLCELL_X8 FILLER_0_34_157 ();
 FILLCELL_X16 FILLER_0_34_170 ();
 FILLCELL_X2 FILLER_0_34_186 ();
 FILLCELL_X2 FILLER_0_34_190 ();
 FILLCELL_X2 FILLER_0_34_194 ();
 FILLCELL_X1 FILLER_0_34_196 ();
 FILLCELL_X4 FILLER_0_34_199 ();
 FILLCELL_X1 FILLER_0_34_203 ();
 FILLCELL_X4 FILLER_0_34_219 ();
 FILLCELL_X2 FILLER_0_34_223 ();
 FILLCELL_X1 FILLER_0_34_225 ();
 FILLCELL_X2 FILLER_0_34_232 ();
 FILLCELL_X4 FILLER_0_34_242 ();
 FILLCELL_X8 FILLER_0_34_255 ();
 FILLCELL_X1 FILLER_0_34_263 ();
 FILLCELL_X2 FILLER_0_34_272 ();
 FILLCELL_X16 FILLER_0_34_276 ();
 FILLCELL_X8 FILLER_0_34_292 ();
 FILLCELL_X2 FILLER_0_34_300 ();
 FILLCELL_X1 FILLER_0_34_302 ();
 FILLCELL_X1 FILLER_0_34_305 ();
 FILLCELL_X2 FILLER_0_34_310 ();
 FILLCELL_X1 FILLER_0_34_312 ();
 FILLCELL_X4 FILLER_0_34_315 ();
 FILLCELL_X1 FILLER_0_34_319 ();
 FILLCELL_X2 FILLER_0_34_324 ();
 FILLCELL_X2 FILLER_0_34_330 ();
 FILLCELL_X1 FILLER_0_34_332 ();
 FILLCELL_X2 FILLER_0_34_335 ();
 FILLCELL_X2 FILLER_0_34_347 ();
 FILLCELL_X1 FILLER_0_34_349 ();
 FILLCELL_X2 FILLER_0_34_365 ();
 FILLCELL_X1 FILLER_0_34_367 ();
 FILLCELL_X4 FILLER_0_34_375 ();
 FILLCELL_X2 FILLER_0_34_379 ();
 FILLCELL_X1 FILLER_0_34_381 ();
 FILLCELL_X1 FILLER_0_34_385 ();
 FILLCELL_X2 FILLER_0_34_393 ();
 FILLCELL_X4 FILLER_0_34_398 ();
 FILLCELL_X8 FILLER_0_34_406 ();
 FILLCELL_X4 FILLER_0_34_414 ();
 FILLCELL_X2 FILLER_0_34_418 ();
 FILLCELL_X1 FILLER_0_34_420 ();
 FILLCELL_X4 FILLER_0_34_424 ();
 FILLCELL_X1 FILLER_0_34_428 ();
 FILLCELL_X4 FILLER_0_34_436 ();
 FILLCELL_X16 FILLER_0_34_448 ();
 FILLCELL_X4 FILLER_0_34_464 ();
 FILLCELL_X2 FILLER_0_35_1 ();
 FILLCELL_X4 FILLER_0_35_6 ();
 FILLCELL_X2 FILLER_0_35_28 ();
 FILLCELL_X16 FILLER_0_35_33 ();
 FILLCELL_X2 FILLER_0_35_52 ();
 FILLCELL_X8 FILLER_0_35_60 ();
 FILLCELL_X4 FILLER_0_35_68 ();
 FILLCELL_X16 FILLER_0_35_77 ();
 FILLCELL_X1 FILLER_0_35_99 ();
 FILLCELL_X1 FILLER_0_35_103 ();
 FILLCELL_X2 FILLER_0_35_107 ();
 FILLCELL_X1 FILLER_0_35_109 ();
 FILLCELL_X16 FILLER_0_35_113 ();
 FILLCELL_X2 FILLER_0_35_129 ();
 FILLCELL_X1 FILLER_0_35_131 ();
 FILLCELL_X4 FILLER_0_35_145 ();
 FILLCELL_X1 FILLER_0_35_149 ();
 FILLCELL_X1 FILLER_0_35_159 ();
 FILLCELL_X2 FILLER_0_35_190 ();
 FILLCELL_X8 FILLER_0_35_198 ();
 FILLCELL_X1 FILLER_0_35_206 ();
 FILLCELL_X2 FILLER_0_35_222 ();
 FILLCELL_X1 FILLER_0_35_224 ();
 FILLCELL_X2 FILLER_0_35_231 ();
 FILLCELL_X1 FILLER_0_35_236 ();
 FILLCELL_X1 FILLER_0_35_247 ();
 FILLCELL_X2 FILLER_0_35_252 ();
 FILLCELL_X1 FILLER_0_35_254 ();
 FILLCELL_X1 FILLER_0_35_262 ();
 FILLCELL_X4 FILLER_0_35_271 ();
 FILLCELL_X2 FILLER_0_35_275 ();
 FILLCELL_X1 FILLER_0_35_277 ();
 FILLCELL_X2 FILLER_0_35_283 ();
 FILLCELL_X1 FILLER_0_35_285 ();
 FILLCELL_X1 FILLER_0_35_288 ();
 FILLCELL_X8 FILLER_0_35_299 ();
 FILLCELL_X2 FILLER_0_35_323 ();
 FILLCELL_X1 FILLER_0_35_339 ();
 FILLCELL_X4 FILLER_0_35_348 ();
 FILLCELL_X2 FILLER_0_35_352 ();
 FILLCELL_X8 FILLER_0_35_360 ();
 FILLCELL_X1 FILLER_0_35_368 ();
 FILLCELL_X4 FILLER_0_35_374 ();
 FILLCELL_X1 FILLER_0_35_378 ();
 FILLCELL_X1 FILLER_0_35_381 ();
 FILLCELL_X1 FILLER_0_35_384 ();
 FILLCELL_X2 FILLER_0_35_389 ();
 FILLCELL_X1 FILLER_0_35_394 ();
 FILLCELL_X4 FILLER_0_35_402 ();
 FILLCELL_X2 FILLER_0_35_406 ();
 FILLCELL_X16 FILLER_0_35_449 ();
 FILLCELL_X2 FILLER_0_35_465 ();
 FILLCELL_X1 FILLER_0_35_467 ();
 FILLCELL_X8 FILLER_0_36_1 ();
 FILLCELL_X4 FILLER_0_36_9 ();
 FILLCELL_X2 FILLER_0_36_52 ();
 FILLCELL_X16 FILLER_0_36_57 ();
 FILLCELL_X1 FILLER_0_36_75 ();
 FILLCELL_X1 FILLER_0_36_107 ();
 FILLCELL_X4 FILLER_0_36_117 ();
 FILLCELL_X2 FILLER_0_36_121 ();
 FILLCELL_X4 FILLER_0_36_139 ();
 FILLCELL_X1 FILLER_0_36_143 ();
 FILLCELL_X2 FILLER_0_36_149 ();
 FILLCELL_X8 FILLER_0_36_176 ();
 FILLCELL_X4 FILLER_0_36_184 ();
 FILLCELL_X2 FILLER_0_36_188 ();
 FILLCELL_X8 FILLER_0_36_198 ();
 FILLCELL_X1 FILLER_0_36_206 ();
 FILLCELL_X4 FILLER_0_36_222 ();
 FILLCELL_X2 FILLER_0_36_226 ();
 FILLCELL_X2 FILLER_0_36_232 ();
 FILLCELL_X4 FILLER_0_36_241 ();
 FILLCELL_X2 FILLER_0_36_251 ();
 FILLCELL_X1 FILLER_0_36_253 ();
 FILLCELL_X4 FILLER_0_36_256 ();
 FILLCELL_X2 FILLER_0_36_260 ();
 FILLCELL_X1 FILLER_0_36_262 ();
 FILLCELL_X1 FILLER_0_36_267 ();
 FILLCELL_X2 FILLER_0_36_277 ();
 FILLCELL_X4 FILLER_0_36_286 ();
 FILLCELL_X1 FILLER_0_36_290 ();
 FILLCELL_X4 FILLER_0_36_298 ();
 FILLCELL_X1 FILLER_0_36_302 ();
 FILLCELL_X1 FILLER_0_36_329 ();
 FILLCELL_X1 FILLER_0_36_333 ();
 FILLCELL_X4 FILLER_0_36_343 ();
 FILLCELL_X1 FILLER_0_36_347 ();
 FILLCELL_X4 FILLER_0_36_358 ();
 FILLCELL_X2 FILLER_0_36_366 ();
 FILLCELL_X1 FILLER_0_36_368 ();
 FILLCELL_X4 FILLER_0_36_389 ();
 FILLCELL_X2 FILLER_0_36_393 ();
 FILLCELL_X1 FILLER_0_36_407 ();
 FILLCELL_X8 FILLER_0_36_414 ();
 FILLCELL_X1 FILLER_0_36_422 ();
 FILLCELL_X2 FILLER_0_36_435 ();
 FILLCELL_X16 FILLER_0_36_445 ();
 FILLCELL_X4 FILLER_0_36_461 ();
 FILLCELL_X2 FILLER_0_36_465 ();
 FILLCELL_X1 FILLER_0_36_467 ();
 FILLCELL_X8 FILLER_0_37_1 ();
 FILLCELL_X4 FILLER_0_37_18 ();
 FILLCELL_X2 FILLER_0_37_22 ();
 FILLCELL_X1 FILLER_0_37_27 ();
 FILLCELL_X1 FILLER_0_37_37 ();
 FILLCELL_X4 FILLER_0_37_40 ();
 FILLCELL_X1 FILLER_0_37_44 ();
 FILLCELL_X16 FILLER_0_37_52 ();
 FILLCELL_X2 FILLER_0_37_68 ();
 FILLCELL_X1 FILLER_0_37_77 ();
 FILLCELL_X1 FILLER_0_37_81 ();
 FILLCELL_X1 FILLER_0_37_84 ();
 FILLCELL_X2 FILLER_0_37_88 ();
 FILLCELL_X2 FILLER_0_37_92 ();
 FILLCELL_X1 FILLER_0_37_94 ();
 FILLCELL_X2 FILLER_0_37_104 ();
 FILLCELL_X16 FILLER_0_37_113 ();
 FILLCELL_X4 FILLER_0_37_129 ();
 FILLCELL_X2 FILLER_0_37_133 ();
 FILLCELL_X1 FILLER_0_37_135 ();
 FILLCELL_X8 FILLER_0_37_153 ();
 FILLCELL_X4 FILLER_0_37_161 ();
 FILLCELL_X2 FILLER_0_37_165 ();
 FILLCELL_X1 FILLER_0_37_173 ();
 FILLCELL_X8 FILLER_0_37_177 ();
 FILLCELL_X4 FILLER_0_37_185 ();
 FILLCELL_X1 FILLER_0_37_189 ();
 FILLCELL_X4 FILLER_0_37_193 ();
 FILLCELL_X1 FILLER_0_37_197 ();
 FILLCELL_X8 FILLER_0_37_200 ();
 FILLCELL_X4 FILLER_0_37_218 ();
 FILLCELL_X1 FILLER_0_37_222 ();
 FILLCELL_X1 FILLER_0_37_227 ();
 FILLCELL_X4 FILLER_0_37_232 ();
 FILLCELL_X2 FILLER_0_37_236 ();
 FILLCELL_X1 FILLER_0_37_238 ();
 FILLCELL_X8 FILLER_0_37_253 ();
 FILLCELL_X1 FILLER_0_37_263 ();
 FILLCELL_X2 FILLER_0_37_271 ();
 FILLCELL_X1 FILLER_0_37_298 ();
 FILLCELL_X16 FILLER_0_37_302 ();
 FILLCELL_X4 FILLER_0_37_318 ();
 FILLCELL_X1 FILLER_0_37_322 ();
 FILLCELL_X2 FILLER_0_37_326 ();
 FILLCELL_X1 FILLER_0_37_331 ();
 FILLCELL_X2 FILLER_0_37_336 ();
 FILLCELL_X1 FILLER_0_37_338 ();
 FILLCELL_X4 FILLER_0_37_347 ();
 FILLCELL_X2 FILLER_0_37_351 ();
 FILLCELL_X1 FILLER_0_37_365 ();
 FILLCELL_X4 FILLER_0_37_379 ();
 FILLCELL_X1 FILLER_0_37_383 ();
 FILLCELL_X4 FILLER_0_37_387 ();
 FILLCELL_X1 FILLER_0_37_391 ();
 FILLCELL_X8 FILLER_0_37_394 ();
 FILLCELL_X4 FILLER_0_37_402 ();
 FILLCELL_X1 FILLER_0_37_420 ();
 FILLCELL_X2 FILLER_0_37_432 ();
 FILLCELL_X16 FILLER_0_37_446 ();
 FILLCELL_X4 FILLER_0_37_462 ();
 FILLCELL_X2 FILLER_0_37_466 ();
 FILLCELL_X1 FILLER_0_38_7 ();
 FILLCELL_X4 FILLER_0_38_20 ();
 FILLCELL_X4 FILLER_0_38_33 ();
 FILLCELL_X1 FILLER_0_38_37 ();
 FILLCELL_X1 FILLER_0_38_41 ();
 FILLCELL_X2 FILLER_0_38_48 ();
 FILLCELL_X1 FILLER_0_38_50 ();
 FILLCELL_X1 FILLER_0_38_62 ();
 FILLCELL_X4 FILLER_0_38_69 ();
 FILLCELL_X1 FILLER_0_38_73 ();
 FILLCELL_X4 FILLER_0_38_76 ();
 FILLCELL_X2 FILLER_0_38_80 ();
 FILLCELL_X1 FILLER_0_38_82 ();
 FILLCELL_X4 FILLER_0_38_93 ();
 FILLCELL_X1 FILLER_0_38_97 ();
 FILLCELL_X4 FILLER_0_38_100 ();
 FILLCELL_X2 FILLER_0_38_104 ();
 FILLCELL_X8 FILLER_0_38_157 ();
 FILLCELL_X2 FILLER_0_38_165 ();
 FILLCELL_X1 FILLER_0_38_167 ();
 FILLCELL_X1 FILLER_0_38_170 ();
 FILLCELL_X1 FILLER_0_38_176 ();
 FILLCELL_X4 FILLER_0_38_187 ();
 FILLCELL_X1 FILLER_0_38_191 ();
 FILLCELL_X1 FILLER_0_38_202 ();
 FILLCELL_X8 FILLER_0_38_205 ();
 FILLCELL_X8 FILLER_0_38_216 ();
 FILLCELL_X2 FILLER_0_38_224 ();
 FILLCELL_X1 FILLER_0_38_232 ();
 FILLCELL_X2 FILLER_0_38_237 ();
 FILLCELL_X4 FILLER_0_38_246 ();
 FILLCELL_X4 FILLER_0_38_259 ();
 FILLCELL_X1 FILLER_0_38_263 ();
 FILLCELL_X2 FILLER_0_38_276 ();
 FILLCELL_X1 FILLER_0_38_281 ();
 FILLCELL_X8 FILLER_0_38_293 ();
 FILLCELL_X4 FILLER_0_38_305 ();
 FILLCELL_X2 FILLER_0_38_316 ();
 FILLCELL_X2 FILLER_0_38_321 ();
 FILLCELL_X2 FILLER_0_38_326 ();
 FILLCELL_X1 FILLER_0_38_331 ();
 FILLCELL_X1 FILLER_0_38_338 ();
 FILLCELL_X8 FILLER_0_38_342 ();
 FILLCELL_X1 FILLER_0_38_350 ();
 FILLCELL_X2 FILLER_0_38_355 ();
 FILLCELL_X8 FILLER_0_38_363 ();
 FILLCELL_X4 FILLER_0_38_374 ();
 FILLCELL_X1 FILLER_0_38_378 ();
 FILLCELL_X2 FILLER_0_38_404 ();
 FILLCELL_X16 FILLER_0_38_440 ();
 FILLCELL_X8 FILLER_0_38_456 ();
 FILLCELL_X4 FILLER_0_38_464 ();
 FILLCELL_X1 FILLER_0_39_4 ();
 FILLCELL_X1 FILLER_0_39_9 ();
 FILLCELL_X1 FILLER_0_39_12 ();
 FILLCELL_X2 FILLER_0_39_17 ();
 FILLCELL_X2 FILLER_0_39_21 ();
 FILLCELL_X1 FILLER_0_39_23 ();
 FILLCELL_X1 FILLER_0_39_30 ();
 FILLCELL_X2 FILLER_0_39_34 ();
 FILLCELL_X4 FILLER_0_39_39 ();
 FILLCELL_X1 FILLER_0_39_43 ();
 FILLCELL_X1 FILLER_0_39_47 ();
 FILLCELL_X8 FILLER_0_39_52 ();
 FILLCELL_X4 FILLER_0_39_66 ();
 FILLCELL_X2 FILLER_0_39_70 ();
 FILLCELL_X1 FILLER_0_39_72 ();
 FILLCELL_X8 FILLER_0_39_80 ();
 FILLCELL_X4 FILLER_0_39_88 ();
 FILLCELL_X1 FILLER_0_39_92 ();
 FILLCELL_X1 FILLER_0_39_96 ();
 FILLCELL_X4 FILLER_0_39_106 ();
 FILLCELL_X2 FILLER_0_39_110 ();
 FILLCELL_X1 FILLER_0_39_112 ();
 FILLCELL_X2 FILLER_0_39_119 ();
 FILLCELL_X16 FILLER_0_39_124 ();
 FILLCELL_X4 FILLER_0_39_150 ();
 FILLCELL_X1 FILLER_0_39_154 ();
 FILLCELL_X2 FILLER_0_39_165 ();
 FILLCELL_X1 FILLER_0_39_167 ();
 FILLCELL_X1 FILLER_0_39_171 ();
 FILLCELL_X8 FILLER_0_39_180 ();
 FILLCELL_X2 FILLER_0_39_188 ();
 FILLCELL_X1 FILLER_0_39_199 ();
 FILLCELL_X4 FILLER_0_39_204 ();
 FILLCELL_X2 FILLER_0_39_208 ();
 FILLCELL_X1 FILLER_0_39_210 ();
 FILLCELL_X2 FILLER_0_39_213 ();
 FILLCELL_X8 FILLER_0_39_228 ();
 FILLCELL_X2 FILLER_0_39_236 ();
 FILLCELL_X16 FILLER_0_39_248 ();
 FILLCELL_X4 FILLER_0_39_264 ();
 FILLCELL_X1 FILLER_0_39_281 ();
 FILLCELL_X4 FILLER_0_39_285 ();
 FILLCELL_X1 FILLER_0_39_289 ();
 FILLCELL_X1 FILLER_0_39_293 ();
 FILLCELL_X8 FILLER_0_39_317 ();
 FILLCELL_X1 FILLER_0_39_325 ();
 FILLCELL_X2 FILLER_0_39_332 ();
 FILLCELL_X1 FILLER_0_39_334 ();
 FILLCELL_X4 FILLER_0_39_338 ();
 FILLCELL_X2 FILLER_0_39_342 ();
 FILLCELL_X2 FILLER_0_39_353 ();
 FILLCELL_X8 FILLER_0_39_358 ();
 FILLCELL_X1 FILLER_0_39_366 ();
 FILLCELL_X4 FILLER_0_39_371 ();
 FILLCELL_X2 FILLER_0_39_378 ();
 FILLCELL_X1 FILLER_0_39_380 ();
 FILLCELL_X2 FILLER_0_39_391 ();
 FILLCELL_X1 FILLER_0_39_393 ();
 FILLCELL_X4 FILLER_0_39_398 ();
 FILLCELL_X2 FILLER_0_39_402 ();
 FILLCELL_X8 FILLER_0_39_412 ();
 FILLCELL_X4 FILLER_0_39_420 ();
 FILLCELL_X2 FILLER_0_39_430 ();
 FILLCELL_X16 FILLER_0_39_448 ();
 FILLCELL_X4 FILLER_0_39_464 ();
 FILLCELL_X1 FILLER_0_40_1 ();
 FILLCELL_X1 FILLER_0_40_18 ();
 FILLCELL_X2 FILLER_0_40_23 ();
 FILLCELL_X1 FILLER_0_40_28 ();
 FILLCELL_X2 FILLER_0_40_32 ();
 FILLCELL_X4 FILLER_0_40_40 ();
 FILLCELL_X2 FILLER_0_40_44 ();
 FILLCELL_X4 FILLER_0_40_52 ();
 FILLCELL_X16 FILLER_0_40_61 ();
 FILLCELL_X4 FILLER_0_40_77 ();
 FILLCELL_X4 FILLER_0_40_93 ();
 FILLCELL_X2 FILLER_0_40_97 ();
 FILLCELL_X1 FILLER_0_40_99 ();
 FILLCELL_X8 FILLER_0_40_107 ();
 FILLCELL_X1 FILLER_0_40_115 ();
 FILLCELL_X4 FILLER_0_40_126 ();
 FILLCELL_X4 FILLER_0_40_138 ();
 FILLCELL_X1 FILLER_0_40_142 ();
 FILLCELL_X2 FILLER_0_40_146 ();
 FILLCELL_X2 FILLER_0_40_158 ();
 FILLCELL_X1 FILLER_0_40_160 ();
 FILLCELL_X2 FILLER_0_40_165 ();
 FILLCELL_X1 FILLER_0_40_167 ();
 FILLCELL_X2 FILLER_0_40_176 ();
 FILLCELL_X1 FILLER_0_40_189 ();
 FILLCELL_X4 FILLER_0_40_193 ();
 FILLCELL_X1 FILLER_0_40_200 ();
 FILLCELL_X1 FILLER_0_40_204 ();
 FILLCELL_X1 FILLER_0_40_208 ();
 FILLCELL_X1 FILLER_0_40_213 ();
 FILLCELL_X8 FILLER_0_40_224 ();
 FILLCELL_X2 FILLER_0_40_232 ();
 FILLCELL_X1 FILLER_0_40_234 ();
 FILLCELL_X2 FILLER_0_40_243 ();
 FILLCELL_X1 FILLER_0_40_248 ();
 FILLCELL_X1 FILLER_0_40_271 ();
 FILLCELL_X1 FILLER_0_40_275 ();
 FILLCELL_X4 FILLER_0_40_289 ();
 FILLCELL_X8 FILLER_0_40_312 ();
 FILLCELL_X2 FILLER_0_40_337 ();
 FILLCELL_X1 FILLER_0_40_350 ();
 FILLCELL_X2 FILLER_0_40_355 ();
 FILLCELL_X2 FILLER_0_40_365 ();
 FILLCELL_X4 FILLER_0_40_389 ();
 FILLCELL_X1 FILLER_0_40_393 ();
 FILLCELL_X2 FILLER_0_40_401 ();
 FILLCELL_X1 FILLER_0_40_403 ();
 FILLCELL_X8 FILLER_0_40_413 ();
 FILLCELL_X2 FILLER_0_40_428 ();
 FILLCELL_X2 FILLER_0_40_436 ();
 FILLCELL_X16 FILLER_0_40_444 ();
 FILLCELL_X8 FILLER_0_40_460 ();
 FILLCELL_X2 FILLER_0_41_1 ();
 FILLCELL_X1 FILLER_0_41_3 ();
 FILLCELL_X4 FILLER_0_41_14 ();
 FILLCELL_X2 FILLER_0_41_18 ();
 FILLCELL_X4 FILLER_0_41_55 ();
 FILLCELL_X1 FILLER_0_41_59 ();
 FILLCELL_X2 FILLER_0_41_67 ();
 FILLCELL_X1 FILLER_0_41_69 ();
 FILLCELL_X2 FILLER_0_41_79 ();
 FILLCELL_X4 FILLER_0_41_93 ();
 FILLCELL_X1 FILLER_0_41_114 ();
 FILLCELL_X1 FILLER_0_41_120 ();
 FILLCELL_X4 FILLER_0_41_125 ();
 FILLCELL_X1 FILLER_0_41_129 ();
 FILLCELL_X8 FILLER_0_41_136 ();
 FILLCELL_X2 FILLER_0_41_144 ();
 FILLCELL_X1 FILLER_0_41_146 ();
 FILLCELL_X4 FILLER_0_41_173 ();
 FILLCELL_X2 FILLER_0_41_177 ();
 FILLCELL_X1 FILLER_0_41_179 ();
 FILLCELL_X1 FILLER_0_41_182 ();
 FILLCELL_X2 FILLER_0_41_194 ();
 FILLCELL_X1 FILLER_0_41_201 ();
 FILLCELL_X2 FILLER_0_41_204 ();
 FILLCELL_X8 FILLER_0_41_212 ();
 FILLCELL_X4 FILLER_0_41_220 ();
 FILLCELL_X2 FILLER_0_41_224 ();
 FILLCELL_X1 FILLER_0_41_226 ();
 FILLCELL_X16 FILLER_0_41_244 ();
 FILLCELL_X1 FILLER_0_41_268 ();
 FILLCELL_X2 FILLER_0_41_273 ();
 FILLCELL_X2 FILLER_0_41_279 ();
 FILLCELL_X2 FILLER_0_41_285 ();
 FILLCELL_X2 FILLER_0_41_295 ();
 FILLCELL_X1 FILLER_0_41_297 ();
 FILLCELL_X8 FILLER_0_41_321 ();
 FILLCELL_X4 FILLER_0_41_329 ();
 FILLCELL_X2 FILLER_0_41_333 ();
 FILLCELL_X1 FILLER_0_41_335 ();
 FILLCELL_X8 FILLER_0_41_355 ();
 FILLCELL_X1 FILLER_0_41_363 ();
 FILLCELL_X8 FILLER_0_41_367 ();
 FILLCELL_X2 FILLER_0_41_378 ();
 FILLCELL_X2 FILLER_0_41_383 ();
 FILLCELL_X4 FILLER_0_41_403 ();
 FILLCELL_X2 FILLER_0_41_407 ();
 FILLCELL_X4 FILLER_0_41_416 ();
 FILLCELL_X2 FILLER_0_41_420 ();
 FILLCELL_X4 FILLER_0_41_430 ();
 FILLCELL_X16 FILLER_0_41_445 ();
 FILLCELL_X4 FILLER_0_41_461 ();
 FILLCELL_X2 FILLER_0_41_465 ();
 FILLCELL_X1 FILLER_0_41_467 ();
 FILLCELL_X1 FILLER_0_42_1 ();
 FILLCELL_X8 FILLER_0_42_28 ();
 FILLCELL_X2 FILLER_0_42_36 ();
 FILLCELL_X1 FILLER_0_42_38 ();
 FILLCELL_X2 FILLER_0_42_44 ();
 FILLCELL_X2 FILLER_0_42_54 ();
 FILLCELL_X1 FILLER_0_42_60 ();
 FILLCELL_X2 FILLER_0_42_78 ();
 FILLCELL_X1 FILLER_0_42_80 ();
 FILLCELL_X8 FILLER_0_42_94 ();
 FILLCELL_X4 FILLER_0_42_105 ();
 FILLCELL_X2 FILLER_0_42_109 ();
 FILLCELL_X1 FILLER_0_42_111 ();
 FILLCELL_X2 FILLER_0_42_120 ();
 FILLCELL_X4 FILLER_0_42_127 ();
 FILLCELL_X4 FILLER_0_42_134 ();
 FILLCELL_X1 FILLER_0_42_138 ();
 FILLCELL_X2 FILLER_0_42_148 ();
 FILLCELL_X4 FILLER_0_42_175 ();
 FILLCELL_X1 FILLER_0_42_185 ();
 FILLCELL_X1 FILLER_0_42_189 ();
 FILLCELL_X4 FILLER_0_42_193 ();
 FILLCELL_X1 FILLER_0_42_197 ();
 FILLCELL_X4 FILLER_0_42_202 ();
 FILLCELL_X2 FILLER_0_42_206 ();
 FILLCELL_X1 FILLER_0_42_208 ();
 FILLCELL_X8 FILLER_0_42_211 ();
 FILLCELL_X4 FILLER_0_42_219 ();
 FILLCELL_X1 FILLER_0_42_223 ();
 FILLCELL_X4 FILLER_0_42_229 ();
 FILLCELL_X2 FILLER_0_42_233 ();
 FILLCELL_X1 FILLER_0_42_235 ();
 FILLCELL_X4 FILLER_0_42_240 ();
 FILLCELL_X2 FILLER_0_42_244 ();
 FILLCELL_X1 FILLER_0_42_246 ();
 FILLCELL_X4 FILLER_0_42_260 ();
 FILLCELL_X1 FILLER_0_42_264 ();
 FILLCELL_X8 FILLER_0_42_269 ();
 FILLCELL_X4 FILLER_0_42_277 ();
 FILLCELL_X1 FILLER_0_42_281 ();
 FILLCELL_X1 FILLER_0_42_293 ();
 FILLCELL_X8 FILLER_0_42_298 ();
 FILLCELL_X4 FILLER_0_42_306 ();
 FILLCELL_X2 FILLER_0_42_310 ();
 FILLCELL_X4 FILLER_0_42_328 ();
 FILLCELL_X2 FILLER_0_42_332 ();
 FILLCELL_X8 FILLER_0_42_337 ();
 FILLCELL_X4 FILLER_0_42_345 ();
 FILLCELL_X2 FILLER_0_42_352 ();
 FILLCELL_X4 FILLER_0_42_367 ();
 FILLCELL_X1 FILLER_0_42_380 ();
 FILLCELL_X2 FILLER_0_42_384 ();
 FILLCELL_X1 FILLER_0_42_386 ();
 FILLCELL_X2 FILLER_0_42_398 ();
 FILLCELL_X1 FILLER_0_42_400 ();
 FILLCELL_X1 FILLER_0_42_405 ();
 FILLCELL_X4 FILLER_0_42_419 ();
 FILLCELL_X2 FILLER_0_42_430 ();
 FILLCELL_X2 FILLER_0_42_435 ();
 FILLCELL_X1 FILLER_0_42_437 ();
 FILLCELL_X16 FILLER_0_42_440 ();
 FILLCELL_X8 FILLER_0_42_456 ();
 FILLCELL_X4 FILLER_0_42_464 ();
 FILLCELL_X8 FILLER_0_43_1 ();
 FILLCELL_X2 FILLER_0_43_9 ();
 FILLCELL_X1 FILLER_0_43_11 ();
 FILLCELL_X1 FILLER_0_43_15 ();
 FILLCELL_X1 FILLER_0_43_21 ();
 FILLCELL_X8 FILLER_0_43_32 ();
 FILLCELL_X4 FILLER_0_43_40 ();
 FILLCELL_X1 FILLER_0_43_44 ();
 FILLCELL_X2 FILLER_0_43_50 ();
 FILLCELL_X1 FILLER_0_43_52 ();
 FILLCELL_X8 FILLER_0_43_62 ();
 FILLCELL_X1 FILLER_0_43_74 ();
 FILLCELL_X8 FILLER_0_43_89 ();
 FILLCELL_X4 FILLER_0_43_97 ();
 FILLCELL_X2 FILLER_0_43_101 ();
 FILLCELL_X2 FILLER_0_43_107 ();
 FILLCELL_X4 FILLER_0_43_113 ();
 FILLCELL_X2 FILLER_0_43_117 ();
 FILLCELL_X1 FILLER_0_43_119 ();
 FILLCELL_X2 FILLER_0_43_124 ();
 FILLCELL_X1 FILLER_0_43_126 ();
 FILLCELL_X1 FILLER_0_43_133 ();
 FILLCELL_X2 FILLER_0_43_151 ();
 FILLCELL_X8 FILLER_0_43_167 ();
 FILLCELL_X2 FILLER_0_43_175 ();
 FILLCELL_X1 FILLER_0_43_177 ();
 FILLCELL_X2 FILLER_0_43_181 ();
 FILLCELL_X1 FILLER_0_43_183 ();
 FILLCELL_X2 FILLER_0_43_196 ();
 FILLCELL_X2 FILLER_0_43_200 ();
 FILLCELL_X1 FILLER_0_43_202 ();
 FILLCELL_X1 FILLER_0_43_223 ();
 FILLCELL_X1 FILLER_0_43_257 ();
 FILLCELL_X4 FILLER_0_43_262 ();
 FILLCELL_X2 FILLER_0_43_270 ();
 FILLCELL_X8 FILLER_0_43_280 ();
 FILLCELL_X4 FILLER_0_43_288 ();
 FILLCELL_X2 FILLER_0_43_311 ();
 FILLCELL_X1 FILLER_0_43_313 ();
 FILLCELL_X2 FILLER_0_43_317 ();
 FILLCELL_X1 FILLER_0_43_338 ();
 FILLCELL_X2 FILLER_0_43_347 ();
 FILLCELL_X2 FILLER_0_43_352 ();
 FILLCELL_X2 FILLER_0_43_357 ();
 FILLCELL_X2 FILLER_0_43_363 ();
 FILLCELL_X1 FILLER_0_43_365 ();
 FILLCELL_X4 FILLER_0_43_371 ();
 FILLCELL_X16 FILLER_0_43_381 ();
 FILLCELL_X8 FILLER_0_43_397 ();
 FILLCELL_X1 FILLER_0_43_405 ();
 FILLCELL_X2 FILLER_0_43_413 ();
 FILLCELL_X4 FILLER_0_43_418 ();
 FILLCELL_X1 FILLER_0_43_422 ();
 FILLCELL_X4 FILLER_0_43_432 ();
 FILLCELL_X1 FILLER_0_43_436 ();
 FILLCELL_X8 FILLER_0_43_454 ();
 FILLCELL_X4 FILLER_0_43_462 ();
 FILLCELL_X2 FILLER_0_43_466 ();
 FILLCELL_X1 FILLER_0_44_4 ();
 FILLCELL_X2 FILLER_0_44_8 ();
 FILLCELL_X2 FILLER_0_44_20 ();
 FILLCELL_X1 FILLER_0_44_22 ();
 FILLCELL_X4 FILLER_0_44_39 ();
 FILLCELL_X2 FILLER_0_44_46 ();
 FILLCELL_X8 FILLER_0_44_55 ();
 FILLCELL_X2 FILLER_0_44_63 ();
 FILLCELL_X2 FILLER_0_44_68 ();
 FILLCELL_X4 FILLER_0_44_73 ();
 FILLCELL_X2 FILLER_0_44_87 ();
 FILLCELL_X1 FILLER_0_44_95 ();
 FILLCELL_X4 FILLER_0_44_98 ();
 FILLCELL_X1 FILLER_0_44_102 ();
 FILLCELL_X8 FILLER_0_44_124 ();
 FILLCELL_X4 FILLER_0_44_147 ();
 FILLCELL_X1 FILLER_0_44_151 ();
 FILLCELL_X16 FILLER_0_44_155 ();
 FILLCELL_X4 FILLER_0_44_171 ();
 FILLCELL_X2 FILLER_0_44_175 ();
 FILLCELL_X4 FILLER_0_44_179 ();
 FILLCELL_X1 FILLER_0_44_183 ();
 FILLCELL_X4 FILLER_0_44_187 ();
 FILLCELL_X2 FILLER_0_44_191 ();
 FILLCELL_X1 FILLER_0_44_193 ();
 FILLCELL_X4 FILLER_0_44_199 ();
 FILLCELL_X1 FILLER_0_44_203 ();
 FILLCELL_X2 FILLER_0_44_207 ();
 FILLCELL_X4 FILLER_0_44_219 ();
 FILLCELL_X2 FILLER_0_44_231 ();
 FILLCELL_X2 FILLER_0_44_256 ();
 FILLCELL_X1 FILLER_0_44_258 ();
 FILLCELL_X1 FILLER_0_44_273 ();
 FILLCELL_X1 FILLER_0_44_278 ();
 FILLCELL_X2 FILLER_0_44_290 ();
 FILLCELL_X4 FILLER_0_44_295 ();
 FILLCELL_X4 FILLER_0_44_303 ();
 FILLCELL_X2 FILLER_0_44_307 ();
 FILLCELL_X1 FILLER_0_44_309 ();
 FILLCELL_X4 FILLER_0_44_317 ();
 FILLCELL_X2 FILLER_0_44_321 ();
 FILLCELL_X1 FILLER_0_44_323 ();
 FILLCELL_X2 FILLER_0_44_328 ();
 FILLCELL_X1 FILLER_0_44_330 ();
 FILLCELL_X2 FILLER_0_44_338 ();
 FILLCELL_X1 FILLER_0_44_340 ();
 FILLCELL_X8 FILLER_0_44_345 ();
 FILLCELL_X1 FILLER_0_44_357 ();
 FILLCELL_X1 FILLER_0_44_362 ();
 FILLCELL_X1 FILLER_0_44_367 ();
 FILLCELL_X4 FILLER_0_44_372 ();
 FILLCELL_X1 FILLER_0_44_376 ();
 FILLCELL_X1 FILLER_0_44_387 ();
 FILLCELL_X4 FILLER_0_44_391 ();
 FILLCELL_X2 FILLER_0_44_395 ();
 FILLCELL_X2 FILLER_0_44_413 ();
 FILLCELL_X1 FILLER_0_44_415 ();
 FILLCELL_X2 FILLER_0_44_423 ();
 FILLCELL_X1 FILLER_0_44_429 ();
 FILLCELL_X2 FILLER_0_44_436 ();
 FILLCELL_X16 FILLER_0_44_444 ();
 FILLCELL_X8 FILLER_0_44_460 ();
 FILLCELL_X4 FILLER_0_45_1 ();
 FILLCELL_X1 FILLER_0_45_5 ();
 FILLCELL_X4 FILLER_0_45_10 ();
 FILLCELL_X1 FILLER_0_45_14 ();
 FILLCELL_X2 FILLER_0_45_24 ();
 FILLCELL_X2 FILLER_0_45_31 ();
 FILLCELL_X2 FILLER_0_45_37 ();
 FILLCELL_X1 FILLER_0_45_39 ();
 FILLCELL_X2 FILLER_0_45_45 ();
 FILLCELL_X1 FILLER_0_45_47 ();
 FILLCELL_X8 FILLER_0_45_53 ();
 FILLCELL_X4 FILLER_0_45_61 ();
 FILLCELL_X2 FILLER_0_45_65 ();
 FILLCELL_X2 FILLER_0_45_74 ();
 FILLCELL_X1 FILLER_0_45_76 ();
 FILLCELL_X2 FILLER_0_45_87 ();
 FILLCELL_X1 FILLER_0_45_94 ();
 FILLCELL_X1 FILLER_0_45_144 ();
 FILLCELL_X16 FILLER_0_45_157 ();
 FILLCELL_X2 FILLER_0_45_173 ();
 FILLCELL_X1 FILLER_0_45_175 ();
 FILLCELL_X2 FILLER_0_45_180 ();
 FILLCELL_X1 FILLER_0_45_182 ();
 FILLCELL_X4 FILLER_0_45_191 ();
 FILLCELL_X2 FILLER_0_45_199 ();
 FILLCELL_X2 FILLER_0_45_204 ();
 FILLCELL_X4 FILLER_0_45_216 ();
 FILLCELL_X2 FILLER_0_45_249 ();
 FILLCELL_X8 FILLER_0_45_284 ();
 FILLCELL_X1 FILLER_0_45_295 ();
 FILLCELL_X8 FILLER_0_45_303 ();
 FILLCELL_X4 FILLER_0_45_311 ();
 FILLCELL_X2 FILLER_0_45_321 ();
 FILLCELL_X1 FILLER_0_45_323 ();
 FILLCELL_X8 FILLER_0_45_336 ();
 FILLCELL_X1 FILLER_0_45_347 ();
 FILLCELL_X2 FILLER_0_45_351 ();
 FILLCELL_X1 FILLER_0_45_353 ();
 FILLCELL_X8 FILLER_0_45_357 ();
 FILLCELL_X4 FILLER_0_45_365 ();
 FILLCELL_X2 FILLER_0_45_369 ();
 FILLCELL_X1 FILLER_0_45_374 ();
 FILLCELL_X2 FILLER_0_45_384 ();
 FILLCELL_X8 FILLER_0_45_392 ();
 FILLCELL_X1 FILLER_0_45_400 ();
 FILLCELL_X16 FILLER_0_45_407 ();
 FILLCELL_X4 FILLER_0_45_423 ();
 FILLCELL_X4 FILLER_0_45_435 ();
 FILLCELL_X2 FILLER_0_45_439 ();
 FILLCELL_X1 FILLER_0_45_441 ();
 FILLCELL_X16 FILLER_0_45_450 ();
 FILLCELL_X2 FILLER_0_45_466 ();
 FILLCELL_X4 FILLER_0_46_1 ();
 FILLCELL_X2 FILLER_0_46_5 ();
 FILLCELL_X1 FILLER_0_46_45 ();
 FILLCELL_X4 FILLER_0_46_49 ();
 FILLCELL_X2 FILLER_0_46_53 ();
 FILLCELL_X1 FILLER_0_46_60 ();
 FILLCELL_X8 FILLER_0_46_63 ();
 FILLCELL_X2 FILLER_0_46_76 ();
 FILLCELL_X8 FILLER_0_46_83 ();
 FILLCELL_X4 FILLER_0_46_91 ();
 FILLCELL_X2 FILLER_0_46_95 ();
 FILLCELL_X1 FILLER_0_46_103 ();
 FILLCELL_X4 FILLER_0_46_118 ();
 FILLCELL_X2 FILLER_0_46_122 ();
 FILLCELL_X2 FILLER_0_46_135 ();
 FILLCELL_X2 FILLER_0_46_140 ();
 FILLCELL_X2 FILLER_0_46_151 ();
 FILLCELL_X2 FILLER_0_46_156 ();
 FILLCELL_X1 FILLER_0_46_158 ();
 FILLCELL_X1 FILLER_0_46_179 ();
 FILLCELL_X2 FILLER_0_46_182 ();
 FILLCELL_X1 FILLER_0_46_184 ();
 FILLCELL_X2 FILLER_0_46_190 ();
 FILLCELL_X2 FILLER_0_46_194 ();
 FILLCELL_X4 FILLER_0_46_199 ();
 FILLCELL_X2 FILLER_0_46_203 ();
 FILLCELL_X1 FILLER_0_46_205 ();
 FILLCELL_X8 FILLER_0_46_209 ();
 FILLCELL_X4 FILLER_0_46_217 ();
 FILLCELL_X2 FILLER_0_46_230 ();
 FILLCELL_X4 FILLER_0_46_236 ();
 FILLCELL_X1 FILLER_0_46_240 ();
 FILLCELL_X2 FILLER_0_46_261 ();
 FILLCELL_X2 FILLER_0_46_274 ();
 FILLCELL_X1 FILLER_0_46_276 ();
 FILLCELL_X1 FILLER_0_46_284 ();
 FILLCELL_X4 FILLER_0_46_291 ();
 FILLCELL_X2 FILLER_0_46_295 ();
 FILLCELL_X4 FILLER_0_46_304 ();
 FILLCELL_X1 FILLER_0_46_308 ();
 FILLCELL_X1 FILLER_0_46_317 ();
 FILLCELL_X4 FILLER_0_46_322 ();
 FILLCELL_X1 FILLER_0_46_326 ();
 FILLCELL_X1 FILLER_0_46_367 ();
 FILLCELL_X4 FILLER_0_46_372 ();
 FILLCELL_X1 FILLER_0_46_376 ();
 FILLCELL_X2 FILLER_0_46_391 ();
 FILLCELL_X1 FILLER_0_46_411 ();
 FILLCELL_X2 FILLER_0_46_416 ();
 FILLCELL_X1 FILLER_0_46_418 ();
 FILLCELL_X1 FILLER_0_46_429 ();
 FILLCELL_X1 FILLER_0_46_433 ();
 FILLCELL_X16 FILLER_0_46_448 ();
 FILLCELL_X4 FILLER_0_46_464 ();
 FILLCELL_X8 FILLER_0_47_4 ();
 FILLCELL_X8 FILLER_0_47_16 ();
 FILLCELL_X4 FILLER_0_47_24 ();
 FILLCELL_X2 FILLER_0_47_28 ();
 FILLCELL_X1 FILLER_0_47_30 ();
 FILLCELL_X1 FILLER_0_47_47 ();
 FILLCELL_X4 FILLER_0_47_54 ();
 FILLCELL_X2 FILLER_0_47_58 ();
 FILLCELL_X8 FILLER_0_47_67 ();
 FILLCELL_X2 FILLER_0_47_75 ();
 FILLCELL_X4 FILLER_0_47_82 ();
 FILLCELL_X1 FILLER_0_47_86 ();
 FILLCELL_X2 FILLER_0_47_105 ();
 FILLCELL_X1 FILLER_0_47_107 ();
 FILLCELL_X8 FILLER_0_47_116 ();
 FILLCELL_X1 FILLER_0_47_124 ();
 FILLCELL_X2 FILLER_0_47_127 ();
 FILLCELL_X1 FILLER_0_47_129 ();
 FILLCELL_X32 FILLER_0_47_132 ();
 FILLCELL_X1 FILLER_0_47_166 ();
 FILLCELL_X1 FILLER_0_47_180 ();
 FILLCELL_X1 FILLER_0_47_204 ();
 FILLCELL_X2 FILLER_0_47_207 ();
 FILLCELL_X8 FILLER_0_47_212 ();
 FILLCELL_X2 FILLER_0_47_220 ();
 FILLCELL_X8 FILLER_0_47_227 ();
 FILLCELL_X4 FILLER_0_47_235 ();
 FILLCELL_X2 FILLER_0_47_239 ();
 FILLCELL_X1 FILLER_0_47_241 ();
 FILLCELL_X1 FILLER_0_47_261 ();
 FILLCELL_X2 FILLER_0_47_269 ();
 FILLCELL_X2 FILLER_0_47_285 ();
 FILLCELL_X8 FILLER_0_47_294 ();
 FILLCELL_X4 FILLER_0_47_302 ();
 FILLCELL_X2 FILLER_0_47_312 ();
 FILLCELL_X1 FILLER_0_47_314 ();
 FILLCELL_X1 FILLER_0_47_319 ();
 FILLCELL_X2 FILLER_0_47_324 ();
 FILLCELL_X1 FILLER_0_47_326 ();
 FILLCELL_X8 FILLER_0_47_330 ();
 FILLCELL_X1 FILLER_0_47_338 ();
 FILLCELL_X1 FILLER_0_47_352 ();
 FILLCELL_X2 FILLER_0_47_365 ();
 FILLCELL_X1 FILLER_0_47_374 ();
 FILLCELL_X2 FILLER_0_47_377 ();
 FILLCELL_X8 FILLER_0_47_383 ();
 FILLCELL_X1 FILLER_0_47_406 ();
 FILLCELL_X2 FILLER_0_47_410 ();
 FILLCELL_X1 FILLER_0_47_412 ();
 FILLCELL_X2 FILLER_0_47_417 ();
 FILLCELL_X1 FILLER_0_47_419 ();
 FILLCELL_X4 FILLER_0_47_430 ();
 FILLCELL_X2 FILLER_0_47_434 ();
 FILLCELL_X1 FILLER_0_47_436 ();
 FILLCELL_X16 FILLER_0_47_448 ();
 FILLCELL_X4 FILLER_0_47_464 ();
 FILLCELL_X32 FILLER_0_48_1 ();
 FILLCELL_X8 FILLER_0_48_33 ();
 FILLCELL_X1 FILLER_0_48_41 ();
 FILLCELL_X16 FILLER_0_48_49 ();
 FILLCELL_X2 FILLER_0_48_65 ();
 FILLCELL_X1 FILLER_0_48_79 ();
 FILLCELL_X8 FILLER_0_48_94 ();
 FILLCELL_X2 FILLER_0_48_102 ();
 FILLCELL_X8 FILLER_0_48_110 ();
 FILLCELL_X4 FILLER_0_48_118 ();
 FILLCELL_X1 FILLER_0_48_135 ();
 FILLCELL_X1 FILLER_0_48_139 ();
 FILLCELL_X2 FILLER_0_48_147 ();
 FILLCELL_X16 FILLER_0_48_152 ();
 FILLCELL_X4 FILLER_0_48_168 ();
 FILLCELL_X2 FILLER_0_48_172 ();
 FILLCELL_X2 FILLER_0_48_178 ();
 FILLCELL_X1 FILLER_0_48_180 ();
 FILLCELL_X1 FILLER_0_48_185 ();
 FILLCELL_X4 FILLER_0_48_215 ();
 FILLCELL_X1 FILLER_0_48_219 ();
 FILLCELL_X4 FILLER_0_48_225 ();
 FILLCELL_X4 FILLER_0_48_234 ();
 FILLCELL_X2 FILLER_0_48_238 ();
 FILLCELL_X1 FILLER_0_48_240 ();
 FILLCELL_X2 FILLER_0_48_246 ();
 FILLCELL_X2 FILLER_0_48_252 ();
 FILLCELL_X1 FILLER_0_48_254 ();
 FILLCELL_X2 FILLER_0_48_264 ();
 FILLCELL_X1 FILLER_0_48_266 ();
 FILLCELL_X8 FILLER_0_48_271 ();
 FILLCELL_X2 FILLER_0_48_283 ();
 FILLCELL_X2 FILLER_0_48_290 ();
 FILLCELL_X1 FILLER_0_48_292 ();
 FILLCELL_X2 FILLER_0_48_301 ();
 FILLCELL_X2 FILLER_0_48_320 ();
 FILLCELL_X1 FILLER_0_48_336 ();
 FILLCELL_X8 FILLER_0_48_343 ();
 FILLCELL_X2 FILLER_0_48_351 ();
 FILLCELL_X1 FILLER_0_48_353 ();
 FILLCELL_X4 FILLER_0_48_367 ();
 FILLCELL_X2 FILLER_0_48_371 ();
 FILLCELL_X1 FILLER_0_48_373 ();
 FILLCELL_X1 FILLER_0_48_377 ();
 FILLCELL_X8 FILLER_0_48_388 ();
 FILLCELL_X4 FILLER_0_48_396 ();
 FILLCELL_X2 FILLER_0_48_400 ();
 FILLCELL_X4 FILLER_0_48_410 ();
 FILLCELL_X2 FILLER_0_48_414 ();
 FILLCELL_X8 FILLER_0_48_423 ();
 FILLCELL_X2 FILLER_0_48_431 ();
 FILLCELL_X1 FILLER_0_48_437 ();
 FILLCELL_X16 FILLER_0_48_441 ();
 FILLCELL_X8 FILLER_0_48_457 ();
 FILLCELL_X2 FILLER_0_48_465 ();
 FILLCELL_X1 FILLER_0_48_467 ();
 FILLCELL_X32 FILLER_0_49_1 ();
 FILLCELL_X32 FILLER_0_49_33 ();
 FILLCELL_X4 FILLER_0_49_65 ();
 FILLCELL_X2 FILLER_0_49_69 ();
 FILLCELL_X1 FILLER_0_49_71 ();
 FILLCELL_X8 FILLER_0_49_77 ();
 FILLCELL_X2 FILLER_0_49_85 ();
 FILLCELL_X4 FILLER_0_49_90 ();
 FILLCELL_X2 FILLER_0_49_94 ();
 FILLCELL_X8 FILLER_0_49_98 ();
 FILLCELL_X1 FILLER_0_49_106 ();
 FILLCELL_X8 FILLER_0_49_112 ();
 FILLCELL_X4 FILLER_0_49_120 ();
 FILLCELL_X8 FILLER_0_49_129 ();
 FILLCELL_X4 FILLER_0_49_137 ();
 FILLCELL_X1 FILLER_0_49_143 ();
 FILLCELL_X1 FILLER_0_49_148 ();
 FILLCELL_X8 FILLER_0_49_158 ();
 FILLCELL_X4 FILLER_0_49_166 ();
 FILLCELL_X1 FILLER_0_49_181 ();
 FILLCELL_X2 FILLER_0_49_185 ();
 FILLCELL_X1 FILLER_0_49_187 ();
 FILLCELL_X2 FILLER_0_49_193 ();
 FILLCELL_X8 FILLER_0_49_203 ();
 FILLCELL_X2 FILLER_0_49_217 ();
 FILLCELL_X1 FILLER_0_49_219 ();
 FILLCELL_X1 FILLER_0_49_248 ();
 FILLCELL_X16 FILLER_0_49_257 ();
 FILLCELL_X2 FILLER_0_49_273 ();
 FILLCELL_X1 FILLER_0_49_275 ();
 FILLCELL_X4 FILLER_0_49_284 ();
 FILLCELL_X1 FILLER_0_49_288 ();
 FILLCELL_X2 FILLER_0_49_292 ();
 FILLCELL_X1 FILLER_0_49_298 ();
 FILLCELL_X2 FILLER_0_49_302 ();
 FILLCELL_X2 FILLER_0_49_307 ();
 FILLCELL_X2 FILLER_0_49_313 ();
 FILLCELL_X8 FILLER_0_49_319 ();
 FILLCELL_X1 FILLER_0_49_327 ();
 FILLCELL_X4 FILLER_0_49_340 ();
 FILLCELL_X2 FILLER_0_49_344 ();
 FILLCELL_X8 FILLER_0_49_366 ();
 FILLCELL_X4 FILLER_0_49_377 ();
 FILLCELL_X2 FILLER_0_49_381 ();
 FILLCELL_X1 FILLER_0_49_386 ();
 FILLCELL_X4 FILLER_0_49_397 ();
 FILLCELL_X2 FILLER_0_49_404 ();
 FILLCELL_X8 FILLER_0_49_417 ();
 FILLCELL_X4 FILLER_0_49_425 ();
 FILLCELL_X2 FILLER_0_49_429 ();
 FILLCELL_X1 FILLER_0_49_431 ();
 FILLCELL_X8 FILLER_0_49_453 ();
 FILLCELL_X4 FILLER_0_49_461 ();
 FILLCELL_X2 FILLER_0_49_465 ();
 FILLCELL_X1 FILLER_0_49_467 ();
 FILLCELL_X32 FILLER_0_50_1 ();
 FILLCELL_X32 FILLER_0_50_33 ();
 FILLCELL_X16 FILLER_0_50_65 ();
 FILLCELL_X4 FILLER_0_50_81 ();
 FILLCELL_X2 FILLER_0_50_85 ();
 FILLCELL_X4 FILLER_0_50_102 ();
 FILLCELL_X2 FILLER_0_50_106 ();
 FILLCELL_X1 FILLER_0_50_108 ();
 FILLCELL_X4 FILLER_0_50_116 ();
 FILLCELL_X2 FILLER_0_50_149 ();
 FILLCELL_X8 FILLER_0_50_160 ();
 FILLCELL_X4 FILLER_0_50_168 ();
 FILLCELL_X2 FILLER_0_50_172 ();
 FILLCELL_X1 FILLER_0_50_174 ();
 FILLCELL_X1 FILLER_0_50_192 ();
 FILLCELL_X1 FILLER_0_50_265 ();
 FILLCELL_X2 FILLER_0_50_282 ();
 FILLCELL_X1 FILLER_0_50_284 ();
 FILLCELL_X4 FILLER_0_50_290 ();
 FILLCELL_X4 FILLER_0_50_300 ();
 FILLCELL_X2 FILLER_0_50_307 ();
 FILLCELL_X4 FILLER_0_50_317 ();
 FILLCELL_X2 FILLER_0_50_321 ();
 FILLCELL_X2 FILLER_0_50_337 ();
 FILLCELL_X2 FILLER_0_50_355 ();
 FILLCELL_X1 FILLER_0_50_357 ();
 FILLCELL_X4 FILLER_0_50_361 ();
 FILLCELL_X4 FILLER_0_50_368 ();
 FILLCELL_X2 FILLER_0_50_372 ();
 FILLCELL_X1 FILLER_0_50_374 ();
 FILLCELL_X2 FILLER_0_50_401 ();
 FILLCELL_X1 FILLER_0_50_414 ();
 FILLCELL_X4 FILLER_0_50_422 ();
 FILLCELL_X2 FILLER_0_50_426 ();
 FILLCELL_X1 FILLER_0_50_443 ();
 FILLCELL_X16 FILLER_0_50_446 ();
 FILLCELL_X4 FILLER_0_50_462 ();
 FILLCELL_X2 FILLER_0_50_466 ();
 FILLCELL_X32 FILLER_0_51_1 ();
 FILLCELL_X32 FILLER_0_51_33 ();
 FILLCELL_X32 FILLER_0_51_65 ();
 FILLCELL_X32 FILLER_0_51_97 ();
 FILLCELL_X2 FILLER_0_51_129 ();
 FILLCELL_X1 FILLER_0_51_131 ();
 FILLCELL_X4 FILLER_0_51_136 ();
 FILLCELL_X1 FILLER_0_51_140 ();
 FILLCELL_X4 FILLER_0_51_155 ();
 FILLCELL_X1 FILLER_0_51_161 ();
 FILLCELL_X1 FILLER_0_51_165 ();
 FILLCELL_X4 FILLER_0_51_168 ();
 FILLCELL_X1 FILLER_0_51_177 ();
 FILLCELL_X1 FILLER_0_51_181 ();
 FILLCELL_X1 FILLER_0_51_225 ();
 FILLCELL_X2 FILLER_0_51_234 ();
 FILLCELL_X2 FILLER_0_51_241 ();
 FILLCELL_X2 FILLER_0_51_247 ();
 FILLCELL_X8 FILLER_0_51_252 ();
 FILLCELL_X4 FILLER_0_51_260 ();
 FILLCELL_X2 FILLER_0_51_264 ();
 FILLCELL_X1 FILLER_0_51_266 ();
 FILLCELL_X1 FILLER_0_51_270 ();
 FILLCELL_X2 FILLER_0_51_275 ();
 FILLCELL_X4 FILLER_0_51_290 ();
 FILLCELL_X2 FILLER_0_51_294 ();
 FILLCELL_X4 FILLER_0_51_298 ();
 FILLCELL_X2 FILLER_0_51_302 ();
 FILLCELL_X1 FILLER_0_51_304 ();
 FILLCELL_X2 FILLER_0_51_307 ();
 FILLCELL_X8 FILLER_0_51_312 ();
 FILLCELL_X2 FILLER_0_51_320 ();
 FILLCELL_X2 FILLER_0_51_331 ();
 FILLCELL_X1 FILLER_0_51_333 ();
 FILLCELL_X2 FILLER_0_51_362 ();
 FILLCELL_X2 FILLER_0_51_372 ();
 FILLCELL_X2 FILLER_0_51_377 ();
 FILLCELL_X4 FILLER_0_51_385 ();
 FILLCELL_X1 FILLER_0_51_389 ();
 FILLCELL_X8 FILLER_0_51_393 ();
 FILLCELL_X2 FILLER_0_51_407 ();
 FILLCELL_X32 FILLER_0_51_435 ();
 FILLCELL_X1 FILLER_0_51_467 ();
 FILLCELL_X32 FILLER_0_52_1 ();
 FILLCELL_X32 FILLER_0_52_33 ();
 FILLCELL_X32 FILLER_0_52_65 ();
 FILLCELL_X16 FILLER_0_52_97 ();
 FILLCELL_X4 FILLER_0_52_113 ();
 FILLCELL_X1 FILLER_0_52_144 ();
 FILLCELL_X1 FILLER_0_52_148 ();
 FILLCELL_X1 FILLER_0_52_157 ();
 FILLCELL_X2 FILLER_0_52_161 ();
 FILLCELL_X2 FILLER_0_52_172 ();
 FILLCELL_X1 FILLER_0_52_174 ();
 FILLCELL_X1 FILLER_0_52_185 ();
 FILLCELL_X1 FILLER_0_52_203 ();
 FILLCELL_X1 FILLER_0_52_217 ();
 FILLCELL_X1 FILLER_0_52_226 ();
 FILLCELL_X1 FILLER_0_52_239 ();
 FILLCELL_X1 FILLER_0_52_243 ();
 FILLCELL_X1 FILLER_0_52_254 ();
 FILLCELL_X2 FILLER_0_52_267 ();
 FILLCELL_X1 FILLER_0_52_269 ();
 FILLCELL_X16 FILLER_0_52_276 ();
 FILLCELL_X1 FILLER_0_52_299 ();
 FILLCELL_X1 FILLER_0_52_308 ();
 FILLCELL_X2 FILLER_0_52_313 ();
 FILLCELL_X8 FILLER_0_52_332 ();
 FILLCELL_X4 FILLER_0_52_340 ();
 FILLCELL_X1 FILLER_0_52_344 ();
 FILLCELL_X4 FILLER_0_52_349 ();
 FILLCELL_X2 FILLER_0_52_353 ();
 FILLCELL_X8 FILLER_0_52_358 ();
 FILLCELL_X1 FILLER_0_52_366 ();
 FILLCELL_X8 FILLER_0_52_371 ();
 FILLCELL_X1 FILLER_0_52_379 ();
 FILLCELL_X4 FILLER_0_52_384 ();
 FILLCELL_X2 FILLER_0_52_388 ();
 FILLCELL_X8 FILLER_0_52_398 ();
 FILLCELL_X2 FILLER_0_52_406 ();
 FILLCELL_X1 FILLER_0_52_408 ();
 FILLCELL_X1 FILLER_0_52_417 ();
 FILLCELL_X1 FILLER_0_52_423 ();
 FILLCELL_X1 FILLER_0_52_426 ();
 FILLCELL_X4 FILLER_0_52_435 ();
 FILLCELL_X2 FILLER_0_52_439 ();
 FILLCELL_X16 FILLER_0_52_450 ();
 FILLCELL_X2 FILLER_0_52_466 ();
 FILLCELL_X32 FILLER_0_53_1 ();
 FILLCELL_X32 FILLER_0_53_33 ();
 FILLCELL_X32 FILLER_0_53_65 ();
 FILLCELL_X16 FILLER_0_53_97 ();
 FILLCELL_X8 FILLER_0_53_113 ();
 FILLCELL_X1 FILLER_0_53_121 ();
 FILLCELL_X1 FILLER_0_53_132 ();
 FILLCELL_X2 FILLER_0_53_135 ();
 FILLCELL_X1 FILLER_0_53_141 ();
 FILLCELL_X1 FILLER_0_53_144 ();
 FILLCELL_X1 FILLER_0_53_148 ();
 FILLCELL_X1 FILLER_0_53_153 ();
 FILLCELL_X4 FILLER_0_53_157 ();
 FILLCELL_X4 FILLER_0_53_164 ();
 FILLCELL_X1 FILLER_0_53_168 ();
 FILLCELL_X1 FILLER_0_53_182 ();
 FILLCELL_X1 FILLER_0_53_211 ();
 FILLCELL_X8 FILLER_0_53_230 ();
 FILLCELL_X2 FILLER_0_53_238 ();
 FILLCELL_X2 FILLER_0_53_243 ();
 FILLCELL_X2 FILLER_0_53_248 ();
 FILLCELL_X2 FILLER_0_53_266 ();
 FILLCELL_X1 FILLER_0_53_268 ();
 FILLCELL_X2 FILLER_0_53_277 ();
 FILLCELL_X1 FILLER_0_53_279 ();
 FILLCELL_X2 FILLER_0_53_290 ();
 FILLCELL_X4 FILLER_0_53_317 ();
 FILLCELL_X2 FILLER_0_53_321 ();
 FILLCELL_X1 FILLER_0_53_331 ();
 FILLCELL_X1 FILLER_0_53_335 ();
 FILLCELL_X1 FILLER_0_53_340 ();
 FILLCELL_X1 FILLER_0_53_345 ();
 FILLCELL_X2 FILLER_0_53_359 ();
 FILLCELL_X4 FILLER_0_53_378 ();
 FILLCELL_X1 FILLER_0_53_382 ();
 FILLCELL_X8 FILLER_0_53_391 ();
 FILLCELL_X2 FILLER_0_53_399 ();
 FILLCELL_X1 FILLER_0_53_401 ();
 FILLCELL_X1 FILLER_0_53_410 ();
 FILLCELL_X8 FILLER_0_53_434 ();
 FILLCELL_X16 FILLER_0_53_451 ();
 FILLCELL_X1 FILLER_0_53_467 ();
 FILLCELL_X32 FILLER_0_54_1 ();
 FILLCELL_X32 FILLER_0_54_33 ();
 FILLCELL_X32 FILLER_0_54_65 ();
 FILLCELL_X16 FILLER_0_54_97 ();
 FILLCELL_X8 FILLER_0_54_113 ();
 FILLCELL_X4 FILLER_0_54_121 ();
 FILLCELL_X1 FILLER_0_54_125 ();
 FILLCELL_X1 FILLER_0_54_148 ();
 FILLCELL_X1 FILLER_0_54_158 ();
 FILLCELL_X2 FILLER_0_54_161 ();
 FILLCELL_X4 FILLER_0_54_166 ();
 FILLCELL_X1 FILLER_0_54_170 ();
 FILLCELL_X1 FILLER_0_54_191 ();
 FILLCELL_X4 FILLER_0_54_241 ();
 FILLCELL_X2 FILLER_0_54_245 ();
 FILLCELL_X2 FILLER_0_54_254 ();
 FILLCELL_X1 FILLER_0_54_256 ();
 FILLCELL_X1 FILLER_0_54_261 ();
 FILLCELL_X4 FILLER_0_54_273 ();
 FILLCELL_X1 FILLER_0_54_280 ();
 FILLCELL_X2 FILLER_0_54_292 ();
 FILLCELL_X1 FILLER_0_54_294 ();
 FILLCELL_X8 FILLER_0_54_298 ();
 FILLCELL_X4 FILLER_0_54_310 ();
 FILLCELL_X1 FILLER_0_54_314 ();
 FILLCELL_X1 FILLER_0_54_319 ();
 FILLCELL_X8 FILLER_0_54_328 ();
 FILLCELL_X1 FILLER_0_54_336 ();
 FILLCELL_X2 FILLER_0_54_344 ();
 FILLCELL_X1 FILLER_0_54_346 ();
 FILLCELL_X2 FILLER_0_54_354 ();
 FILLCELL_X1 FILLER_0_54_359 ();
 FILLCELL_X4 FILLER_0_54_370 ();
 FILLCELL_X4 FILLER_0_54_377 ();
 FILLCELL_X2 FILLER_0_54_381 ();
 FILLCELL_X1 FILLER_0_54_383 ();
 FILLCELL_X1 FILLER_0_54_419 ();
 FILLCELL_X2 FILLER_0_54_423 ();
 FILLCELL_X8 FILLER_0_54_456 ();
 FILLCELL_X4 FILLER_0_54_464 ();
 FILLCELL_X32 FILLER_0_55_1 ();
 FILLCELL_X32 FILLER_0_55_33 ();
 FILLCELL_X32 FILLER_0_55_65 ();
 FILLCELL_X16 FILLER_0_55_97 ();
 FILLCELL_X8 FILLER_0_55_113 ();
 FILLCELL_X4 FILLER_0_55_121 ();
 FILLCELL_X1 FILLER_0_55_133 ();
 FILLCELL_X2 FILLER_0_55_138 ();
 FILLCELL_X1 FILLER_0_55_140 ();
 FILLCELL_X1 FILLER_0_55_146 ();
 FILLCELL_X4 FILLER_0_55_150 ();
 FILLCELL_X1 FILLER_0_55_154 ();
 FILLCELL_X4 FILLER_0_55_161 ();
 FILLCELL_X2 FILLER_0_55_165 ();
 FILLCELL_X1 FILLER_0_55_167 ();
 FILLCELL_X8 FILLER_0_55_238 ();
 FILLCELL_X4 FILLER_0_55_246 ();
 FILLCELL_X1 FILLER_0_55_250 ();
 FILLCELL_X2 FILLER_0_55_254 ();
 FILLCELL_X1 FILLER_0_55_256 ();
 FILLCELL_X4 FILLER_0_55_261 ();
 FILLCELL_X1 FILLER_0_55_265 ();
 FILLCELL_X2 FILLER_0_55_272 ();
 FILLCELL_X1 FILLER_0_55_274 ();
 FILLCELL_X4 FILLER_0_55_283 ();
 FILLCELL_X1 FILLER_0_55_287 ();
 FILLCELL_X1 FILLER_0_55_291 ();
 FILLCELL_X2 FILLER_0_55_298 ();
 FILLCELL_X1 FILLER_0_55_300 ();
 FILLCELL_X1 FILLER_0_55_304 ();
 FILLCELL_X4 FILLER_0_55_319 ();
 FILLCELL_X1 FILLER_0_55_323 ();
 FILLCELL_X2 FILLER_0_55_330 ();
 FILLCELL_X2 FILLER_0_55_335 ();
 FILLCELL_X1 FILLER_0_55_341 ();
 FILLCELL_X1 FILLER_0_55_346 ();
 FILLCELL_X4 FILLER_0_55_354 ();
 FILLCELL_X1 FILLER_0_55_358 ();
 FILLCELL_X8 FILLER_0_55_366 ();
 FILLCELL_X1 FILLER_0_55_374 ();
 FILLCELL_X4 FILLER_0_55_387 ();
 FILLCELL_X1 FILLER_0_55_391 ();
 FILLCELL_X1 FILLER_0_55_399 ();
 FILLCELL_X1 FILLER_0_55_404 ();
 FILLCELL_X1 FILLER_0_55_408 ();
 FILLCELL_X1 FILLER_0_55_413 ();
 FILLCELL_X16 FILLER_0_55_422 ();
 FILLCELL_X8 FILLER_0_55_438 ();
 FILLCELL_X16 FILLER_0_55_448 ();
 FILLCELL_X4 FILLER_0_55_464 ();
 FILLCELL_X32 FILLER_0_56_1 ();
 FILLCELL_X32 FILLER_0_56_33 ();
 FILLCELL_X32 FILLER_0_56_65 ();
 FILLCELL_X16 FILLER_0_56_97 ();
 FILLCELL_X8 FILLER_0_56_113 ();
 FILLCELL_X1 FILLER_0_56_121 ();
 FILLCELL_X1 FILLER_0_56_142 ();
 FILLCELL_X1 FILLER_0_56_148 ();
 FILLCELL_X1 FILLER_0_56_152 ();
 FILLCELL_X2 FILLER_0_56_155 ();
 FILLCELL_X2 FILLER_0_56_161 ();
 FILLCELL_X2 FILLER_0_56_165 ();
 FILLCELL_X1 FILLER_0_56_170 ();
 FILLCELL_X4 FILLER_0_56_177 ();
 FILLCELL_X2 FILLER_0_56_181 ();
 FILLCELL_X4 FILLER_0_56_187 ();
 FILLCELL_X1 FILLER_0_56_200 ();
 FILLCELL_X1 FILLER_0_56_226 ();
 FILLCELL_X4 FILLER_0_56_236 ();
 FILLCELL_X16 FILLER_0_56_251 ();
 FILLCELL_X8 FILLER_0_56_267 ();
 FILLCELL_X4 FILLER_0_56_275 ();
 FILLCELL_X2 FILLER_0_56_279 ();
 FILLCELL_X1 FILLER_0_56_281 ();
 FILLCELL_X1 FILLER_0_56_289 ();
 FILLCELL_X4 FILLER_0_56_303 ();
 FILLCELL_X4 FILLER_0_56_314 ();
 FILLCELL_X1 FILLER_0_56_318 ();
 FILLCELL_X2 FILLER_0_56_331 ();
 FILLCELL_X1 FILLER_0_56_336 ();
 FILLCELL_X1 FILLER_0_56_354 ();
 FILLCELL_X8 FILLER_0_56_358 ();
 FILLCELL_X2 FILLER_0_56_379 ();
 FILLCELL_X4 FILLER_0_56_387 ();
 FILLCELL_X1 FILLER_0_56_391 ();
 FILLCELL_X1 FILLER_0_56_395 ();
 FILLCELL_X2 FILLER_0_56_406 ();
 FILLCELL_X1 FILLER_0_56_408 ();
 FILLCELL_X32 FILLER_0_56_413 ();
 FILLCELL_X16 FILLER_0_56_445 ();
 FILLCELL_X4 FILLER_0_56_461 ();
 FILLCELL_X2 FILLER_0_56_465 ();
 FILLCELL_X1 FILLER_0_56_467 ();
 FILLCELL_X32 FILLER_0_57_1 ();
 FILLCELL_X32 FILLER_0_57_33 ();
 FILLCELL_X32 FILLER_0_57_65 ();
 FILLCELL_X32 FILLER_0_57_97 ();
 FILLCELL_X16 FILLER_0_57_129 ();
 FILLCELL_X2 FILLER_0_57_145 ();
 FILLCELL_X1 FILLER_0_57_147 ();
 FILLCELL_X2 FILLER_0_57_154 ();
 FILLCELL_X1 FILLER_0_57_179 ();
 FILLCELL_X1 FILLER_0_57_222 ();
 FILLCELL_X1 FILLER_0_57_227 ();
 FILLCELL_X1 FILLER_0_57_231 ();
 FILLCELL_X2 FILLER_0_57_250 ();
 FILLCELL_X1 FILLER_0_57_257 ();
 FILLCELL_X2 FILLER_0_57_262 ();
 FILLCELL_X8 FILLER_0_57_275 ();
 FILLCELL_X2 FILLER_0_57_283 ();
 FILLCELL_X8 FILLER_0_57_303 ();
 FILLCELL_X4 FILLER_0_57_311 ();
 FILLCELL_X4 FILLER_0_57_319 ();
 FILLCELL_X2 FILLER_0_57_323 ();
 FILLCELL_X16 FILLER_0_57_331 ();
 FILLCELL_X8 FILLER_0_57_352 ();
 FILLCELL_X4 FILLER_0_57_360 ();
 FILLCELL_X2 FILLER_0_57_364 ();
 FILLCELL_X8 FILLER_0_57_371 ();
 FILLCELL_X1 FILLER_0_57_379 ();
 FILLCELL_X4 FILLER_0_57_383 ();
 FILLCELL_X1 FILLER_0_57_387 ();
 FILLCELL_X32 FILLER_0_57_394 ();
 FILLCELL_X32 FILLER_0_57_426 ();
 FILLCELL_X8 FILLER_0_57_458 ();
 FILLCELL_X2 FILLER_0_57_466 ();
 FILLCELL_X32 FILLER_0_58_1 ();
 FILLCELL_X32 FILLER_0_58_33 ();
 FILLCELL_X32 FILLER_0_58_65 ();
 FILLCELL_X32 FILLER_0_58_97 ();
 FILLCELL_X8 FILLER_0_58_129 ();
 FILLCELL_X4 FILLER_0_58_137 ();
 FILLCELL_X2 FILLER_0_58_144 ();
 FILLCELL_X2 FILLER_0_58_159 ();
 FILLCELL_X1 FILLER_0_58_161 ();
 FILLCELL_X1 FILLER_0_58_165 ();
 FILLCELL_X4 FILLER_0_58_172 ();
 FILLCELL_X2 FILLER_0_58_176 ();
 FILLCELL_X1 FILLER_0_58_178 ();
 FILLCELL_X4 FILLER_0_58_181 ();
 FILLCELL_X1 FILLER_0_58_185 ();
 FILLCELL_X1 FILLER_0_58_195 ();
 FILLCELL_X4 FILLER_0_58_199 ();
 FILLCELL_X1 FILLER_0_58_203 ();
 FILLCELL_X4 FILLER_0_58_211 ();
 FILLCELL_X1 FILLER_0_58_215 ();
 FILLCELL_X1 FILLER_0_58_246 ();
 FILLCELL_X16 FILLER_0_58_271 ();
 FILLCELL_X8 FILLER_0_58_287 ();
 FILLCELL_X1 FILLER_0_58_304 ();
 FILLCELL_X4 FILLER_0_58_310 ();
 FILLCELL_X1 FILLER_0_58_314 ();
 FILLCELL_X4 FILLER_0_58_322 ();
 FILLCELL_X2 FILLER_0_58_326 ();
 FILLCELL_X1 FILLER_0_58_335 ();
 FILLCELL_X8 FILLER_0_58_346 ();
 FILLCELL_X16 FILLER_0_58_357 ();
 FILLCELL_X1 FILLER_0_58_373 ();
 FILLCELL_X32 FILLER_0_58_392 ();
 FILLCELL_X32 FILLER_0_58_424 ();
 FILLCELL_X8 FILLER_0_58_456 ();
 FILLCELL_X4 FILLER_0_58_464 ();
 FILLCELL_X32 FILLER_0_59_1 ();
 FILLCELL_X32 FILLER_0_59_33 ();
 FILLCELL_X32 FILLER_0_59_65 ();
 FILLCELL_X32 FILLER_0_59_97 ();
 FILLCELL_X8 FILLER_0_59_129 ();
 FILLCELL_X4 FILLER_0_59_137 ();
 FILLCELL_X2 FILLER_0_59_141 ();
 FILLCELL_X1 FILLER_0_59_143 ();
 FILLCELL_X1 FILLER_0_59_150 ();
 FILLCELL_X4 FILLER_0_59_155 ();
 FILLCELL_X1 FILLER_0_59_159 ();
 FILLCELL_X2 FILLER_0_59_166 ();
 FILLCELL_X1 FILLER_0_59_168 ();
 FILLCELL_X4 FILLER_0_59_190 ();
 FILLCELL_X8 FILLER_0_59_197 ();
 FILLCELL_X2 FILLER_0_59_205 ();
 FILLCELL_X1 FILLER_0_59_209 ();
 FILLCELL_X1 FILLER_0_59_214 ();
 FILLCELL_X1 FILLER_0_59_223 ();
 FILLCELL_X2 FILLER_0_59_234 ();
 FILLCELL_X1 FILLER_0_59_236 ();
 FILLCELL_X1 FILLER_0_59_240 ();
 FILLCELL_X4 FILLER_0_59_247 ();
 FILLCELL_X2 FILLER_0_59_251 ();
 FILLCELL_X1 FILLER_0_59_255 ();
 FILLCELL_X8 FILLER_0_59_266 ();
 FILLCELL_X1 FILLER_0_59_274 ();
 FILLCELL_X2 FILLER_0_59_277 ();
 FILLCELL_X1 FILLER_0_59_284 ();
 FILLCELL_X1 FILLER_0_59_289 ();
 FILLCELL_X1 FILLER_0_59_295 ();
 FILLCELL_X1 FILLER_0_59_299 ();
 FILLCELL_X2 FILLER_0_59_304 ();
 FILLCELL_X2 FILLER_0_59_314 ();
 FILLCELL_X1 FILLER_0_59_316 ();
 FILLCELL_X1 FILLER_0_59_342 ();
 FILLCELL_X8 FILLER_0_59_364 ();
 FILLCELL_X2 FILLER_0_59_372 ();
 FILLCELL_X32 FILLER_0_59_392 ();
 FILLCELL_X32 FILLER_0_59_424 ();
 FILLCELL_X8 FILLER_0_59_456 ();
 FILLCELL_X4 FILLER_0_59_464 ();
 FILLCELL_X32 FILLER_0_60_1 ();
 FILLCELL_X32 FILLER_0_60_33 ();
 FILLCELL_X32 FILLER_0_60_65 ();
 FILLCELL_X32 FILLER_0_60_97 ();
 FILLCELL_X16 FILLER_0_60_129 ();
 FILLCELL_X2 FILLER_0_60_145 ();
 FILLCELL_X4 FILLER_0_60_149 ();
 FILLCELL_X2 FILLER_0_60_153 ();
 FILLCELL_X16 FILLER_0_60_158 ();
 FILLCELL_X8 FILLER_0_60_182 ();
 FILLCELL_X1 FILLER_0_60_190 ();
 FILLCELL_X1 FILLER_0_60_200 ();
 FILLCELL_X8 FILLER_0_60_214 ();
 FILLCELL_X2 FILLER_0_60_222 ();
 FILLCELL_X1 FILLER_0_60_229 ();
 FILLCELL_X4 FILLER_0_60_235 ();
 FILLCELL_X2 FILLER_0_60_239 ();
 FILLCELL_X2 FILLER_0_60_246 ();
 FILLCELL_X1 FILLER_0_60_248 ();
 FILLCELL_X4 FILLER_0_60_252 ();
 FILLCELL_X4 FILLER_0_60_260 ();
 FILLCELL_X2 FILLER_0_60_264 ();
 FILLCELL_X1 FILLER_0_60_266 ();
 FILLCELL_X8 FILLER_0_60_281 ();
 FILLCELL_X4 FILLER_0_60_289 ();
 FILLCELL_X1 FILLER_0_60_293 ();
 FILLCELL_X8 FILLER_0_60_297 ();
 FILLCELL_X4 FILLER_0_60_305 ();
 FILLCELL_X2 FILLER_0_60_309 ();
 FILLCELL_X1 FILLER_0_60_311 ();
 FILLCELL_X4 FILLER_0_60_315 ();
 FILLCELL_X4 FILLER_0_60_337 ();
 FILLCELL_X2 FILLER_0_60_341 ();
 FILLCELL_X4 FILLER_0_60_348 ();
 FILLCELL_X1 FILLER_0_60_352 ();
 FILLCELL_X1 FILLER_0_60_357 ();
 FILLCELL_X1 FILLER_0_60_367 ();
 FILLCELL_X32 FILLER_0_60_380 ();
 FILLCELL_X32 FILLER_0_60_412 ();
 FILLCELL_X16 FILLER_0_60_444 ();
 FILLCELL_X8 FILLER_0_60_460 ();
 FILLCELL_X32 FILLER_0_61_1 ();
 FILLCELL_X32 FILLER_0_61_33 ();
 FILLCELL_X32 FILLER_0_61_65 ();
 FILLCELL_X32 FILLER_0_61_97 ();
 FILLCELL_X8 FILLER_0_61_129 ();
 FILLCELL_X4 FILLER_0_61_137 ();
 FILLCELL_X1 FILLER_0_61_141 ();
 FILLCELL_X1 FILLER_0_61_145 ();
 FILLCELL_X4 FILLER_0_61_167 ();
 FILLCELL_X1 FILLER_0_61_171 ();
 FILLCELL_X2 FILLER_0_61_188 ();
 FILLCELL_X2 FILLER_0_61_196 ();
 FILLCELL_X1 FILLER_0_61_213 ();
 FILLCELL_X2 FILLER_0_61_220 ();
 FILLCELL_X1 FILLER_0_61_222 ();
 FILLCELL_X8 FILLER_0_61_229 ();
 FILLCELL_X4 FILLER_0_61_237 ();
 FILLCELL_X2 FILLER_0_61_241 ();
 FILLCELL_X16 FILLER_0_61_253 ();
 FILLCELL_X2 FILLER_0_61_269 ();
 FILLCELL_X1 FILLER_0_61_271 ();
 FILLCELL_X2 FILLER_0_61_275 ();
 FILLCELL_X4 FILLER_0_61_284 ();
 FILLCELL_X2 FILLER_0_61_288 ();
 FILLCELL_X1 FILLER_0_61_293 ();
 FILLCELL_X2 FILLER_0_61_300 ();
 FILLCELL_X1 FILLER_0_61_302 ();
 FILLCELL_X1 FILLER_0_61_312 ();
 FILLCELL_X1 FILLER_0_61_331 ();
 FILLCELL_X1 FILLER_0_61_335 ();
 FILLCELL_X1 FILLER_0_61_342 ();
 FILLCELL_X1 FILLER_0_61_352 ();
 FILLCELL_X4 FILLER_0_61_368 ();
 FILLCELL_X2 FILLER_0_61_375 ();
 FILLCELL_X1 FILLER_0_61_377 ();
 FILLCELL_X32 FILLER_0_61_381 ();
 FILLCELL_X32 FILLER_0_61_413 ();
 FILLCELL_X16 FILLER_0_61_445 ();
 FILLCELL_X4 FILLER_0_61_461 ();
 FILLCELL_X2 FILLER_0_61_465 ();
 FILLCELL_X1 FILLER_0_61_467 ();
 FILLCELL_X32 FILLER_0_62_1 ();
 FILLCELL_X32 FILLER_0_62_33 ();
 FILLCELL_X32 FILLER_0_62_65 ();
 FILLCELL_X32 FILLER_0_62_97 ();
 FILLCELL_X8 FILLER_0_62_129 ();
 FILLCELL_X4 FILLER_0_62_137 ();
 FILLCELL_X2 FILLER_0_62_144 ();
 FILLCELL_X8 FILLER_0_62_152 ();
 FILLCELL_X4 FILLER_0_62_160 ();
 FILLCELL_X2 FILLER_0_62_164 ();
 FILLCELL_X1 FILLER_0_62_166 ();
 FILLCELL_X8 FILLER_0_62_170 ();
 FILLCELL_X4 FILLER_0_62_178 ();
 FILLCELL_X2 FILLER_0_62_182 ();
 FILLCELL_X1 FILLER_0_62_184 ();
 FILLCELL_X2 FILLER_0_62_194 ();
 FILLCELL_X16 FILLER_0_62_199 ();
 FILLCELL_X1 FILLER_0_62_215 ();
 FILLCELL_X8 FILLER_0_62_228 ();
 FILLCELL_X4 FILLER_0_62_236 ();
 FILLCELL_X2 FILLER_0_62_240 ();
 FILLCELL_X1 FILLER_0_62_242 ();
 FILLCELL_X16 FILLER_0_62_255 ();
 FILLCELL_X4 FILLER_0_62_271 ();
 FILLCELL_X2 FILLER_0_62_275 ();
 FILLCELL_X2 FILLER_0_62_286 ();
 FILLCELL_X1 FILLER_0_62_288 ();
 FILLCELL_X1 FILLER_0_62_298 ();
 FILLCELL_X1 FILLER_0_62_305 ();
 FILLCELL_X2 FILLER_0_62_315 ();
 FILLCELL_X1 FILLER_0_62_317 ();
 FILLCELL_X2 FILLER_0_62_327 ();
 FILLCELL_X1 FILLER_0_62_338 ();
 FILLCELL_X1 FILLER_0_62_342 ();
 FILLCELL_X1 FILLER_0_62_358 ();
 FILLCELL_X1 FILLER_0_62_368 ();
 FILLCELL_X16 FILLER_0_62_372 ();
 FILLCELL_X32 FILLER_0_62_391 ();
 FILLCELL_X32 FILLER_0_62_423 ();
 FILLCELL_X8 FILLER_0_62_455 ();
 FILLCELL_X4 FILLER_0_62_463 ();
 FILLCELL_X1 FILLER_0_62_467 ();
endmodule
