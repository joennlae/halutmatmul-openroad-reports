module halut_decoder__2864165611389228789 (clk_i,
    decoder_i,
    rst_ni,
    valid_o,
    we_i,
    c_addr_i,
    k_addr_i,
    result_o,
    waddr_i,
    wdata_i);
 input clk_i;
 input decoder_i;
 input rst_ni;
 output valid_o;
 input we_i;
 input [4:0] c_addr_i;
 input [3:0] k_addr_i;
 output [31:0] result_o;
 input [8:0] waddr_i;
 input [7:0] wdata_i;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire net55;
 wire _00534_;
 wire net52;
 wire net51;
 wire _00537_;
 wire net49;
 wire net48;
 wire _00540_;
 wire net46;
 wire net45;
 wire _00543_;
 wire net43;
 wire net42;
 wire _00546_;
 wire net40;
 wire net39;
 wire _00549_;
 wire net37;
 wire net36;
 wire _00552_;
 wire net34;
 wire net33;
 wire _00555_;
 wire net31;
 wire net30;
 wire _00558_;
 wire net28;
 wire net27;
 wire _00561_;
 wire net25;
 wire net24;
 wire _00564_;
 wire net22;
 wire net21;
 wire _00567_;
 wire net19;
 wire net18;
 wire _00570_;
 wire net16;
 wire net15;
 wire _00573_;
 wire net13;
 wire net12;
 wire _00576_;
 wire net10;
 wire net9;
 wire _00579_;
 wire net7;
 wire net6;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire net5;
 wire _00586_;
 wire net4;
 wire _00588_;
 wire _00589_;
 wire net3;
 wire net2;
 wire _00592_;
 wire net1;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ;
 wire _00655_;
 wire _00656_;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ;
 wire _00660_;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire \clknet_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ;
 wire _00686_;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire \clknet_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ;
 wire _00703_;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ;
 wire _00705_;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire \clknet_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ;
 wire clknet_level_2_1_8140__00537_;
 wire clknet_level_1_1_8139__00537_;
 wire clknet_level_0_1_8138__00537_;
 wire clknet_level_2_1_7137__00537_;
 wire clknet_level_1_1_7136__00537_;
 wire clknet_level_0_1_7135__00537_;
 wire clknet_level_2_1_6134__00537_;
 wire clknet_level_1_1_6133__00537_;
 wire clknet_level_0_1_6132__00537_;
 wire clknet_level_2_1_5131__00537_;
 wire clknet_level_1_1_5130__00537_;
 wire clknet_level_0_1_5129__00537_;
 wire clknet_level_2_1_4128__00537_;
 wire clknet_level_1_1_4127__00537_;
 wire clknet_level_0_1_4126__00537_;
 wire clknet_level_2_1_3125__00537_;
 wire clknet_level_1_1_3124__00537_;
 wire clknet_level_0_1_3123__00537_;
 wire clknet_level_2_1_2122__00537_;
 wire clknet_level_1_1_2121__00537_;
 wire clknet_level_0_1_2120__00537_;
 wire clknet_level_2_1_1119__00537_;
 wire clknet_level_1_1_1118__00537_;
 wire clknet_level_0_1_1117__00537_;
 wire clknet_3_7__leaf__00537_;
 wire clknet_3_6__leaf__00537_;
 wire clknet_3_5__leaf__00537_;
 wire clknet_3_4__leaf__00537_;
 wire _00760_;
 wire _00761_;
 wire clknet_3_3__leaf__00537_;
 wire clknet_3_2__leaf__00537_;
 wire clknet_3_1__leaf__00537_;
 wire _00765_;
 wire _00766_;
 wire clknet_3_0__leaf__00537_;
 wire clknet_0__00537_;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ;
 wire _00770_;
 wire _00771_;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ;
 wire _00773_;
 wire \clknet_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ;
 wire _00777_;
 wire \clknet_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ;
 wire _00781_;
 wire \clknet_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ;
 wire _00785_;
 wire \clknet_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire \clknet_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ;
 wire _00795_;
 wire \clknet_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ;
 wire _00799_;
 wire \clknet_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ;
 wire _00803_;
 wire \clknet_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ;
 wire _00807_;
 wire _00808_;
 wire \clknet_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ;
 wire _00812_;
 wire \clknet_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ;
 wire _00816_;
 wire \clknet_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ;
 wire _00820_;
 wire \clknet_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ;
 wire _00830_;
 wire _00831_;
 wire \clknet_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire \clknet_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ;
 wire _00911_;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ;
 wire _00914_;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ;
 wire _00916_;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ;
 wire _00918_;
 wire \clknet_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ;
 wire _00926_;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ;
 wire _00933_;
 wire _00934_;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ;
 wire _00937_;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ;
 wire _00939_;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire \clknet_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ;
 wire _00946_;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ;
 wire _00948_;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ;
 wire _00950_;
 wire \clknet_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ;
 wire _00956_;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ;
 wire _00959_;
 wire _00960_;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ;
 wire _00962_;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ;
 wire _00964_;
 wire \clknet_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ;
 wire _00970_;
 wire _00971_;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ;
 wire _00974_;
 wire _00975_;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire \clknet_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ;
 wire _00989_;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ;
 wire _00996_;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ;
 wire _00998_;
 wire _00999_;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ;
 wire _01002_;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ;
 wire _01004_;
 wire _01005_;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ;
 wire _01007_;
 wire \clknet_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ;
 wire _01009_;
 wire clknet_level_2_1_8242__00534_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire clknet_level_1_1_8241__00534_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire clknet_level_0_1_8240__00534_;
 wire _01021_;
 wire clknet_level_2_1_7239__00534_;
 wire _01023_;
 wire _01024_;
 wire clknet_level_1_1_7238__00534_;
 wire _01026_;
 wire _01027_;
 wire clknet_level_0_1_7237__00534_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire clknet_level_2_1_6236__00534_;
 wire _01034_;
 wire clknet_level_1_1_6235__00534_;
 wire clknet_level_0_1_6234__00534_;
 wire _01037_;
 wire _01038_;
 wire clknet_level_2_1_5233__00534_;
 wire clknet_level_1_1_5232__00534_;
 wire clknet_level_0_1_5231__00534_;
 wire _01042_;
 wire clknet_level_2_1_4230__00534_;
 wire clknet_level_1_1_4229__00534_;
 wire _01045_;
 wire _01046_;
 wire clknet_level_0_1_4228__00534_;
 wire clknet_level_2_1_3227__00534_;
 wire clknet_level_1_1_3226__00534_;
 wire _01050_;
 wire clknet_level_0_1_3225__00534_;
 wire clknet_level_2_1_2224__00534_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire clknet_level_1_1_2223__00534_;
 wire _01059_;
 wire clknet_level_0_1_2222__00534_;
 wire clknet_level_2_1_1221__00534_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire clknet_level_1_1_1220__00534_;
 wire clknet_level_0_1_1219__00534_;
 wire clknet_3_7__leaf__00534_;
 wire _01068_;
 wire clknet_3_6__leaf__00534_;
 wire clknet_3_5__leaf__00534_;
 wire clknet_3_4__leaf__00534_;
 wire clknet_3_3__leaf__00534_;
 wire clknet_3_2__leaf__00534_;
 wire clknet_3_1__leaf__00534_;
 wire _01075_;
 wire _01076_;
 wire clknet_3_0__leaf__00534_;
 wire clknet_0__00534_;
 wire clknet_level_5_1_4320__00532_;
 wire clknet_level_4_1_4319__00532_;
 wire _01081_;
 wire clknet_level_3_1_4318__00532_;
 wire clknet_level_2_1_4317__00532_;
 wire _01084_;
 wire clknet_level_1_1_4316__00532_;
 wire clknet_level_0_1_4315__00532_;
 wire clknet_level_5_1_3218__00532_;
 wire clknet_level_4_1_3217__00532_;
 wire clknet_level_3_1_3216__00532_;
 wire clknet_level_2_1_3215__00532_;
 wire _01091_;
 wire clknet_level_1_1_3214__00532_;
 wire clknet_level_0_1_3213__00532_;
 wire clknet_level_5_1_2116__00532_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire clknet_level_4_1_2115__00532_;
 wire clknet_level_3_1_2114__00532_;
 wire clknet_level_2_1_2113__00532_;
 wire _01101_;
 wire _01102_;
 wire clknet_level_1_1_2112__00532_;
 wire clknet_level_0_1_2111__00532_;
 wire clknet_level_5_1_114__00532_;
 wire clknet_level_4_1_113__00532_;
 wire clknet_level_3_1_112__00532_;
 wire clknet_level_2_1_111__00532_;
 wire _01109_;
 wire clknet_level_1_1_110__00532_;
 wire clknet_level_0_1_19__00532_;
 wire clknet_2_3__leaf__00532_;
 wire _01113_;
 wire clknet_2_2__leaf__00532_;
 wire clknet_2_1__leaf__00532_;
 wire clknet_2_0__leaf__00532_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire clknet_0__00532_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire clknet_level_8_1_8479_clk_i;
 wire _01125_;
 wire clknet_level_7_1_8478_clk_i;
 wire clknet_level_6_1_8477_clk_i;
 wire clknet_level_5_1_8476_clk_i;
 wire clknet_level_4_1_8475_clk_i;
 wire clknet_level_3_1_8474_clk_i;
 wire _01131_;
 wire clknet_level_2_1_8473_clk_i;
 wire clknet_level_1_1_8472_clk_i;
 wire _01134_;
 wire clknet_level_0_1_8471_clk_i;
 wire clknet_level_8_1_7470_clk_i;
 wire clknet_level_7_1_7469_clk_i;
 wire clknet_level_6_1_7468_clk_i;
 wire _01139_;
 wire _01140_;
 wire clknet_level_5_1_7467_clk_i;
 wire clknet_level_4_1_7466_clk_i;
 wire _01143_;
 wire _01144_;
 wire clknet_level_3_1_7465_clk_i;
 wire clknet_level_2_1_7464_clk_i;
 wire clknet_level_1_1_7463_clk_i;
 wire _01148_;
 wire _01149_;
 wire clknet_level_0_1_7462_clk_i;
 wire clknet_level_8_1_6461_clk_i;
 wire clknet_level_7_1_6460_clk_i;
 wire clknet_level_6_1_6459_clk_i;
 wire clknet_level_5_1_6458_clk_i;
 wire _01155_;
 wire clknet_level_4_1_6457_clk_i;
 wire clknet_level_3_1_6456_clk_i;
 wire clknet_level_2_1_6455_clk_i;
 wire clknet_level_1_1_6454_clk_i;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire clknet_level_0_1_6453_clk_i;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire clknet_level_8_1_5452_clk_i;
 wire clknet_level_7_1_5451_clk_i;
 wire clknet_level_6_1_5450_clk_i;
 wire _01174_;
 wire clknet_level_5_1_5449_clk_i;
 wire clknet_level_4_1_5448_clk_i;
 wire _01177_;
 wire _01178_;
 wire clknet_level_3_1_5447_clk_i;
 wire _01180_;
 wire _01181_;
 wire clknet_level_2_1_5446_clk_i;
 wire _01183_;
 wire _01184_;
 wire clknet_level_1_1_5445_clk_i;
 wire clknet_level_0_1_5444_clk_i;
 wire clknet_level_8_1_4443_clk_i;
 wire clknet_level_7_1_4442_clk_i;
 wire clknet_level_6_1_4441_clk_i;
 wire _01190_;
 wire clknet_level_5_1_4440_clk_i;
 wire clknet_level_4_1_4439_clk_i;
 wire clknet_level_3_1_4438_clk_i;
 wire _01194_;
 wire _01195_;
 wire clknet_level_2_1_4437_clk_i;
 wire _01197_;
 wire clknet_level_1_1_4436_clk_i;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire clknet_level_0_1_4435_clk_i;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire clknet_level_8_1_3434_clk_i;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire clknet_level_7_1_3433_clk_i;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire clknet_level_6_1_3432_clk_i;
 wire clknet_level_5_1_3431_clk_i;
 wire _01225_;
 wire clknet_level_4_1_3430_clk_i;
 wire clknet_level_3_1_3429_clk_i;
 wire clknet_level_2_1_3428_clk_i;
 wire clknet_level_1_1_3427_clk_i;
 wire clknet_level_0_1_3426_clk_i;
 wire _01231_;
 wire clknet_level_8_1_2425_clk_i;
 wire clknet_level_7_1_2424_clk_i;
 wire clknet_level_6_1_2423_clk_i;
 wire clknet_level_5_1_2422_clk_i;
 wire _01236_;
 wire clknet_level_4_1_2421_clk_i;
 wire clknet_level_3_1_2420_clk_i;
 wire clknet_level_2_1_2419_clk_i;
 wire _01240_;
 wire _01241_;
 wire clknet_level_1_1_2418_clk_i;
 wire clknet_level_0_1_2417_clk_i;
 wire clknet_level_8_1_18_clk_i;
 wire clknet_level_7_1_17_clk_i;
 wire _01246_;
 wire clknet_level_6_1_16_clk_i;
 wire clknet_level_5_1_15_clk_i;
 wire clknet_level_4_1_14_clk_i;
 wire _01250_;
 wire clknet_level_3_1_13_clk_i;
 wire clknet_level_2_1_12_clk_i;
 wire clknet_level_1_1_11_clk_i;
 wire clknet_level_0_1_10_clk_i;
 wire _01255_;
 wire clknet_3_7__leaf_clk_i;
 wire clknet_3_6__leaf_clk_i;
 wire clknet_3_5__leaf_clk_i;
 wire _01259_;
 wire _01260_;
 wire clknet_3_4__leaf_clk_i;
 wire clknet_3_3__leaf_clk_i;
 wire _01263_;
 wire clknet_3_2__leaf_clk_i;
 wire clknet_3_1__leaf_clk_i;
 wire clknet_3_0__leaf_clk_i;
 wire clknet_0_clk_i;
 wire _01268_;
 wire net321;
 wire net320;
 wire net319;
 wire net318;
 wire _01273_;
 wire net317;
 wire _01275_;
 wire _01276_;
 wire net316;
 wire net315;
 wire net314;
 wire _01280_;
 wire net313;
 wire net312;
 wire net311;
 wire _01284_;
 wire net310;
 wire net309;
 wire net308;
 wire _01288_;
 wire net307;
 wire net306;
 wire net305;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire net304;
 wire net303;
 wire _01298_;
 wire _01299_;
 wire net302;
 wire _01301_;
 wire net301;
 wire _01303_;
 wire net300;
 wire _01305_;
 wire net299;
 wire net298;
 wire net297;
 wire _01309_;
 wire _01310_;
 wire net296;
 wire _01312_;
 wire net295;
 wire net294;
 wire _01315_;
 wire net293;
 wire net292;
 wire net291;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire net290;
 wire _01323_;
 wire net289;
 wire net288;
 wire _01326_;
 wire net287;
 wire net286;
 wire net285;
 wire _01330_;
 wire net284;
 wire net283;
 wire _01333_;
 wire _01334_;
 wire net282;
 wire net281;
 wire net280;
 wire net279;
 wire _01339_;
 wire net278;
 wire net277;
 wire _01342_;
 wire net276;
 wire _01344_;
 wire net275;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire net274;
 wire net273;
 wire net272;
 wire net271;
 wire _01356_;
 wire net270;
 wire _01358_;
 wire net269;
 wire _01360_;
 wire net268;
 wire net267;
 wire _01363_;
 wire _01364_;
 wire net266;
 wire _01366_;
 wire net265;
 wire net264;
 wire net263;
 wire _01370_;
 wire net262;
 wire _01372_;
 wire net261;
 wire _01374_;
 wire net260;
 wire _01376_;
 wire _01377_;
 wire net259;
 wire net258;
 wire _01380_;
 wire net257;
 wire _01382_;
 wire net256;
 wire net255;
 wire _01385_;
 wire net254;
 wire _01387_;
 wire _01388_;
 wire net253;
 wire net252;
 wire _01391_;
 wire net251;
 wire net250;
 wire _01394_;
 wire net249;
 wire _01396_;
 wire net248;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire net247;
 wire net246;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire net245;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire net244;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire net243;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire net242;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire net241;
 wire _01437_;
 wire net240;
 wire net239;
 wire _01440_;
 wire net238;
 wire net237;
 wire _01443_;
 wire _01444_;
 wire net236;
 wire _01446_;
 wire net235;
 wire _01448_;
 wire net234;
 wire net233;
 wire net232;
 wire _01452_;
 wire net231;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire net230;
 wire _01463_;
 wire net229;
 wire _01465_;
 wire net228;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire net227;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire net226;
 wire net225;
 wire _01479_;
 wire _01480_;
 wire net224;
 wire _01482_;
 wire net223;
 wire net222;
 wire net221;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire net220;
 wire _01491_;
 wire _01492_;
 wire net219;
 wire net218;
 wire net217;
 wire net216;
 wire _01497_;
 wire net215;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire net214;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire net213;
 wire _01511_;
 wire net212;
 wire _01513_;
 wire _01514_;
 wire net211;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire net210;
 wire net209;
 wire _01521_;
 wire net208;
 wire net207;
 wire _01524_;
 wire net206;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire net205;
 wire net204;
 wire _01531_;
 wire net203;
 wire _01533_;
 wire net202;
 wire net201;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire net200;
 wire _01541_;
 wire _01542_;
 wire net199;
 wire _01544_;
 wire net198;
 wire _01546_;
 wire net197;
 wire net196;
 wire net195;
 wire net194;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire net193;
 wire net192;
 wire _01557_;
 wire net191;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire net190;
 wire _01563_;
 wire net189;
 wire _01565_;
 wire net188;
 wire net187;
 wire _01568_;
 wire net186;
 wire net185;
 wire _01571_;
 wire _01572_;
 wire net184;
 wire _01574_;
 wire net183;
 wire _01576_;
 wire net182;
 wire _01578_;
 wire net181;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire net180;
 wire _01586_;
 wire net179;
 wire net178;
 wire _01589_;
 wire net177;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire net176;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire net175;
 wire _01600_;
 wire _01601_;
 wire net174;
 wire net173;
 wire _01604_;
 wire net172;
 wire _01606_;
 wire net171;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire net170;
 wire net169;
 wire _01613_;
 wire net168;
 wire net167;
 wire _01616_;
 wire _01617_;
 wire net166;
 wire net165;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire net164;
 wire _01625_;
 wire _01626_;
 wire net163;
 wire net162;
 wire _01629_;
 wire net161;
 wire _01631_;
 wire net160;
 wire _01633_;
 wire net159;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire net158;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire net157;
 wire net156;
 wire _01655_;
 wire net155;
 wire _01657_;
 wire net154;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire net153;
 wire net152;
 wire _01666_;
 wire _01667_;
 wire net151;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire net150;
 wire _01673_;
 wire _01674_;
 wire net149;
 wire _01676_;
 wire net148;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire net147;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire net146;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire net145;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire net144;
 wire _01718_;
 wire net143;
 wire net142;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire net141;
 wire _01725_;
 wire net140;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire net139;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire net138;
 wire _01740_;
 wire net137;
 wire _01742_;
 wire net136;
 wire _01744_;
 wire net135;
 wire net134;
 wire _01747_;
 wire _01748_;
 wire net133;
 wire _01750_;
 wire _01751_;
 wire net132;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire net131;
 wire _01757_;
 wire net130;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire net129;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire net128;
 wire net127;
 wire net126;
 wire _01772_;
 wire net125;
 wire net124;
 wire _01775_;
 wire net123;
 wire net122;
 wire _01778_;
 wire net121;
 wire net120;
 wire _01781_;
 wire _01782_;
 wire net119;
 wire net118;
 wire _01785_;
 wire net117;
 wire _01787_;
 wire net116;
 wire net115;
 wire _01790_;
 wire net114;
 wire net113;
 wire _01793_;
 wire _01794_;
 wire net112;
 wire net111;
 wire _01797_;
 wire net110;
 wire net109;
 wire net108;
 wire _01801_;
 wire net107;
 wire _01803_;
 wire net106;
 wire _01805_;
 wire _01806_;
 wire net105;
 wire net104;
 wire _01809_;
 wire net103;
 wire _01811_;
 wire _01812_;
 wire net102;
 wire net101;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire net100;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire net99;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire net98;
 wire _01833_;
 wire _01834_;
 wire net97;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire net96;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire net95;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire net94;
 wire _01854_;
 wire _01855_;
 wire net93;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire net92;
 wire _01864_;
 wire _01865_;
 wire net91;
 wire _01867_;
 wire net90;
 wire _01869_;
 wire net89;
 wire _01871_;
 wire net88;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire net87;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire net86;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire net85;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire net84;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire net83;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire net82;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire net81;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire net80;
 wire _01942_;
 wire net79;
 wire _01944_;
 wire _01945_;
 wire net78;
 wire _01947_;
 wire _01948_;
 wire net77;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire net76;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire net75;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire net74;
 wire _01984_;
 wire _01985_;
 wire net73;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire net72;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire net71;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire net70;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire net69;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire net68;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire net67;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire net66;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire net65;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire net64;
 wire _02348_;
 wire _02349_;
 wire net63;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire net62;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire net61;
 wire _02362_;
 wire _02363_;
 wire net60;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire net59;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire net58;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire net57;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire net56;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire \caddr_n[0] ;
 wire \caddr_n[1] ;
 wire \caddr_n[2] ;
 wire \caddr_n[3] ;
 wire \caddr_n[4] ;
 wire \caddr_q[0] ;
 wire \caddr_q[1] ;
 wire \caddr_q[2] ;
 wire \caddr_q[3] ;
 wire \caddr_q[4] ;
 wire \genblk1.gen_int_accumulation.int_adder.int_long_i[0] ;
 wire \genblk1.gen_int_accumulation.int_adder.int_long_i[10] ;
 wire \genblk1.gen_int_accumulation.int_adder.int_long_i[11] ;
 wire \genblk1.gen_int_accumulation.int_adder.int_long_i[12] ;
 wire \genblk1.gen_int_accumulation.int_adder.int_long_i[13] ;
 wire \genblk1.gen_int_accumulation.int_adder.int_long_i[14] ;
 wire \genblk1.gen_int_accumulation.int_adder.int_long_i[15] ;
 wire \genblk1.gen_int_accumulation.int_adder.int_long_i[16] ;
 wire \genblk1.gen_int_accumulation.int_adder.int_long_i[17] ;
 wire \genblk1.gen_int_accumulation.int_adder.int_long_i[18] ;
 wire \genblk1.gen_int_accumulation.int_adder.int_long_i[19] ;
 wire \genblk1.gen_int_accumulation.int_adder.int_long_i[1] ;
 wire \genblk1.gen_int_accumulation.int_adder.int_long_i[20] ;
 wire \genblk1.gen_int_accumulation.int_adder.int_long_i[21] ;
 wire \genblk1.gen_int_accumulation.int_adder.int_long_i[22] ;
 wire \genblk1.gen_int_accumulation.int_adder.int_long_i[23] ;
 wire \genblk1.gen_int_accumulation.int_adder.int_long_i[24] ;
 wire \genblk1.gen_int_accumulation.int_adder.int_long_i[25] ;
 wire \genblk1.gen_int_accumulation.int_adder.int_long_i[26] ;
 wire \genblk1.gen_int_accumulation.int_adder.int_long_i[27] ;
 wire \genblk1.gen_int_accumulation.int_adder.int_long_i[28] ;
 wire \genblk1.gen_int_accumulation.int_adder.int_long_i[29] ;
 wire \genblk1.gen_int_accumulation.int_adder.int_long_i[2] ;
 wire \genblk1.gen_int_accumulation.int_adder.int_long_i[30] ;
 wire \genblk1.gen_int_accumulation.int_adder.int_long_i[31] ;
 wire \genblk1.gen_int_accumulation.int_adder.int_long_i[3] ;
 wire \genblk1.gen_int_accumulation.int_adder.int_long_i[4] ;
 wire \genblk1.gen_int_accumulation.int_adder.int_long_i[5] ;
 wire \genblk1.gen_int_accumulation.int_adder.int_long_i[6] ;
 wire \genblk1.gen_int_accumulation.int_adder.int_long_i[7] ;
 wire \genblk1.gen_int_accumulation.int_adder.int_long_i[8] ;
 wire \genblk1.gen_int_accumulation.int_adder.int_long_i[9] ;
 wire \genblk1.gen_int_accumulation.int_adder.int_short_converted[0] ;
 wire \genblk1.gen_int_accumulation.int_adder.int_short_converted[10] ;
 wire \genblk1.gen_int_accumulation.int_adder.int_short_converted[1] ;
 wire \genblk1.gen_int_accumulation.int_adder.int_short_converted[2] ;
 wire \genblk1.gen_int_accumulation.int_adder.int_short_converted[3] ;
 wire \genblk1.gen_int_accumulation.int_adder.int_short_converted[4] ;
 wire \genblk1.gen_int_accumulation.int_adder.int_short_converted[5] ;
 wire \genblk1.gen_int_accumulation.int_adder.int_short_converted[6] ;
 wire \lut.cg_we_global.clk_en ;
 wire net54;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.cg_we_global.clk_en ;
 wire net8;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.cg_we_global.en_i ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__0.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__1.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__10.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__11.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__12.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__13.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__14.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__15.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__16.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__17.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__18.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__19.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__2.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__20.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__21.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__22.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__23.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__24.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__25.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__26.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__27.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__28.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__29.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__3.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__30.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__31.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__4.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__5.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__6.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__7.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__8.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__9.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[0][0] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[0][1] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[0][2] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[0][3] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[0][4] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[0][5] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[0][6] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[0][7] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[10][0] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[10][1] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[10][2] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[10][3] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[10][4] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[10][5] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[10][6] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[10][7] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[11][0] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[11][1] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[11][2] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[11][3] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[11][4] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[11][5] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[11][6] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[11][7] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[12][0] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[12][1] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[12][2] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[12][3] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[12][4] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[12][5] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[12][6] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[12][7] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[13][0] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[13][1] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[13][2] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[13][3] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[13][4] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[13][5] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[13][6] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[13][7] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[14][0] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[14][1] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[14][2] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[14][3] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[14][4] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[14][5] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[14][6] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[14][7] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[15][0] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[15][1] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[15][2] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[15][3] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[15][4] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[15][5] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[15][6] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[15][7] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[16][0] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[16][1] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[16][2] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[16][3] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[16][4] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[16][5] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[16][6] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[16][7] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[17][0] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[17][1] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[17][2] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[17][3] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[17][4] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[17][5] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[17][6] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[17][7] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[18][0] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[18][1] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[18][2] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[18][3] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[18][4] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[18][5] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[18][6] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[18][7] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[19][0] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[19][1] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[19][2] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[19][3] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[19][4] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[19][5] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[19][6] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[19][7] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[1][0] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[1][1] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[1][2] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[1][3] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[1][4] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[1][5] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[1][6] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[1][7] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[20][0] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[20][1] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[20][2] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[20][3] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[20][4] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[20][5] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[20][6] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[20][7] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[21][0] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[21][1] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[21][2] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[21][3] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[21][4] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[21][5] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[21][6] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[21][7] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[22][0] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[22][1] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[22][2] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[22][3] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[22][4] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[22][5] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[22][6] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[22][7] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[23][0] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[23][1] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[23][2] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[23][3] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[23][4] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[23][5] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[23][6] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[23][7] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[24][0] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[24][1] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[24][2] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[24][3] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[24][4] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[24][5] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[24][6] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[24][7] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[25][0] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[25][1] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[25][2] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[25][3] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[25][4] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[25][5] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[25][6] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[25][7] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[26][0] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[26][1] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[26][2] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[26][3] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[26][4] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[26][5] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[26][6] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[26][7] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[27][0] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[27][1] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[27][2] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[27][3] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[27][4] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[27][5] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[27][6] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[27][7] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[28][0] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[28][1] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[28][2] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[28][3] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[28][4] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[28][5] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[28][6] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[28][7] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[29][0] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[29][1] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[29][2] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[29][3] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[29][4] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[29][5] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[29][6] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[29][7] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[2][0] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[2][1] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[2][2] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[2][3] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[2][4] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[2][5] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[2][6] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[2][7] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[30][0] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[30][1] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[30][2] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[30][3] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[30][4] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[30][5] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[30][6] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[30][7] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[31][0] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[31][1] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[31][2] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[31][3] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[31][4] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[31][5] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[31][6] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[31][7] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[3][0] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[3][1] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[3][2] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[3][3] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[3][4] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[3][5] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[3][6] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[3][7] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[4][0] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[4][1] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[4][2] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[4][3] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[4][4] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[4][5] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[4][6] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[4][7] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[5][0] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[5][1] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[5][2] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[5][3] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[5][4] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[5][5] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[5][6] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[5][7] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[6][0] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[6][1] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[6][2] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[6][3] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[6][4] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[6][5] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[6][6] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[6][7] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[7][0] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[7][1] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[7][2] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[7][3] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[7][4] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[7][5] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[7][6] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[7][7] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[8][0] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[8][1] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[8][2] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[8][3] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[8][4] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[8][5] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[8][6] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[8][7] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[9][0] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[9][1] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[9][2] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[9][3] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[9][4] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[9][5] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[9][6] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.mem[9][7] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[0] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[1] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[2] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[3] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[4] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[5] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[6] ;
 wire \lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[7] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.cg_we_global.clk_en ;
 wire net11;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.cg_we_global.en_i ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__0.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__1.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__10.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__11.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__12.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__13.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__14.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__15.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__16.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__17.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__18.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__19.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__2.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__20.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__21.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__22.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__23.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__24.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__25.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__26.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__27.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__28.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__29.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__3.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__30.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__31.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__4.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__5.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__6.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__7.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__8.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__9.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[0][0] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[0][1] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[0][2] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[0][3] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[0][4] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[0][5] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[0][6] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[0][7] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[10][0] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[10][1] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[10][2] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[10][3] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[10][4] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[10][5] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[10][6] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[10][7] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[11][0] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[11][1] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[11][2] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[11][3] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[11][4] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[11][5] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[11][6] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[11][7] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[12][0] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[12][1] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[12][2] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[12][3] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[12][4] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[12][5] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[12][6] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[12][7] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[13][0] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[13][1] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[13][2] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[13][3] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[13][4] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[13][5] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[13][6] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[13][7] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[14][0] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[14][1] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[14][2] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[14][3] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[14][4] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[14][5] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[14][6] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[14][7] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[15][0] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[15][1] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[15][2] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[15][3] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[15][4] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[15][5] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[15][6] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[15][7] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[16][0] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[16][1] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[16][2] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[16][3] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[16][4] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[16][5] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[16][6] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[16][7] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[17][0] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[17][1] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[17][2] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[17][3] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[17][4] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[17][5] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[17][6] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[17][7] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[18][0] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[18][1] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[18][2] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[18][3] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[18][4] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[18][5] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[18][6] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[18][7] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[19][0] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[19][1] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[19][2] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[19][3] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[19][4] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[19][5] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[19][6] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[19][7] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[1][0] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[1][1] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[1][2] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[1][3] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[1][4] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[1][5] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[1][6] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[1][7] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[20][0] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[20][1] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[20][2] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[20][3] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[20][4] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[20][5] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[20][6] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[20][7] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[21][0] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[21][1] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[21][2] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[21][3] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[21][4] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[21][5] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[21][6] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[21][7] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[22][0] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[22][1] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[22][2] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[22][3] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[22][4] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[22][5] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[22][6] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[22][7] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[23][0] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[23][1] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[23][2] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[23][3] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[23][4] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[23][5] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[23][6] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[23][7] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[24][0] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[24][1] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[24][2] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[24][3] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[24][4] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[24][5] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[24][6] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[24][7] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[25][0] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[25][1] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[25][2] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[25][3] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[25][4] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[25][5] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[25][6] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[25][7] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[26][0] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[26][1] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[26][2] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[26][3] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[26][4] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[26][5] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[26][6] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[26][7] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[27][0] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[27][1] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[27][2] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[27][3] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[27][4] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[27][5] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[27][6] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[27][7] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[28][0] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[28][1] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[28][2] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[28][3] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[28][4] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[28][5] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[28][6] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[28][7] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[29][0] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[29][1] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[29][2] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[29][3] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[29][4] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[29][5] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[29][6] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[29][7] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[2][0] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[2][1] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[2][2] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[2][3] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[2][4] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[2][5] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[2][6] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[2][7] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[30][0] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[30][1] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[30][2] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[30][3] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[30][4] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[30][5] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[30][6] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[30][7] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[31][0] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[31][1] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[31][2] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[31][3] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[31][4] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[31][5] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[31][6] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[31][7] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[3][0] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[3][1] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[3][2] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[3][3] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[3][4] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[3][5] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[3][6] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[3][7] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[4][0] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[4][1] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[4][2] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[4][3] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[4][4] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[4][5] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[4][6] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[4][7] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[5][0] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[5][1] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[5][2] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[5][3] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[5][4] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[5][5] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[5][6] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[5][7] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[6][0] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[6][1] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[6][2] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[6][3] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[6][4] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[6][5] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[6][6] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[6][7] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[7][0] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[7][1] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[7][2] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[7][3] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[7][4] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[7][5] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[7][6] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[7][7] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[8][0] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[8][1] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[8][2] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[8][3] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[8][4] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[8][5] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[8][6] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[8][7] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[9][0] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[9][1] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[9][2] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[9][3] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[9][4] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[9][5] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[9][6] ;
 wire \lut.gen_sub_units_scm.__1.sub_unit_i.mem[9][7] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.cg_we_global.clk_en ;
 wire net38;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.cg_we_global.en_i ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__0.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__1.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__10.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__11.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__12.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__13.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__14.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__15.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__16.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__17.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__18.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__19.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__2.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__20.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__21.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__22.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__23.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__24.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__25.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__26.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__27.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__28.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__29.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__3.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__30.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__31.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__4.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__5.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__6.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__7.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__8.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__9.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[0][0] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[0][1] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[0][2] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[0][3] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[0][4] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[0][5] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[0][6] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[0][7] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[10][0] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[10][1] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[10][2] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[10][3] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[10][4] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[10][5] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[10][6] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[10][7] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[11][0] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[11][1] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[11][2] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[11][3] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[11][4] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[11][5] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[11][6] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[11][7] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[12][0] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[12][1] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[12][2] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[12][3] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[12][4] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[12][5] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[12][6] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[12][7] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[13][0] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[13][1] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[13][2] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[13][3] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[13][4] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[13][5] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[13][6] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[13][7] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[14][0] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[14][1] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[14][2] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[14][3] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[14][4] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[14][5] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[14][6] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[14][7] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[15][0] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[15][1] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[15][2] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[15][3] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[15][4] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[15][5] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[15][6] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[15][7] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[16][0] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[16][1] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[16][2] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[16][3] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[16][4] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[16][5] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[16][6] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[16][7] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[17][0] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[17][1] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[17][2] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[17][3] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[17][4] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[17][5] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[17][6] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[17][7] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[18][0] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[18][1] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[18][2] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[18][3] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[18][4] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[18][5] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[18][6] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[18][7] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[19][0] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[19][1] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[19][2] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[19][3] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[19][4] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[19][5] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[19][6] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[19][7] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[1][0] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[1][1] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[1][2] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[1][3] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[1][4] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[1][5] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[1][6] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[1][7] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[20][0] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[20][1] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[20][2] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[20][3] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[20][4] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[20][5] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[20][6] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[20][7] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[21][0] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[21][1] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[21][2] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[21][3] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[21][4] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[21][5] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[21][6] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[21][7] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[22][0] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[22][1] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[22][2] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[22][3] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[22][4] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[22][5] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[22][6] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[22][7] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[23][0] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[23][1] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[23][2] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[23][3] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[23][4] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[23][5] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[23][6] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[23][7] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[24][0] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[24][1] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[24][2] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[24][3] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[24][4] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[24][5] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[24][6] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[24][7] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[25][0] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[25][1] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[25][2] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[25][3] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[25][4] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[25][5] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[25][6] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[25][7] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[26][0] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[26][1] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[26][2] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[26][3] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[26][4] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[26][5] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[26][6] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[26][7] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[27][0] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[27][1] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[27][2] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[27][3] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[27][4] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[27][5] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[27][6] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[27][7] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[28][0] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[28][1] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[28][2] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[28][3] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[28][4] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[28][5] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[28][6] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[28][7] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[29][0] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[29][1] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[29][2] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[29][3] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[29][4] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[29][5] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[29][6] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[29][7] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[2][0] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[2][1] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[2][2] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[2][3] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[2][4] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[2][5] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[2][6] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[2][7] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[30][0] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[30][1] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[30][2] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[30][3] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[30][4] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[30][5] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[30][6] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[30][7] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[31][0] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[31][1] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[31][2] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[31][3] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[31][4] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[31][5] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[31][6] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[31][7] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[3][0] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[3][1] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[3][2] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[3][3] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[3][4] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[3][5] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[3][6] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[3][7] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[4][0] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[4][1] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[4][2] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[4][3] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[4][4] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[4][5] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[4][6] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[4][7] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[5][0] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[5][1] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[5][2] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[5][3] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[5][4] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[5][5] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[5][6] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[5][7] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[6][0] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[6][1] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[6][2] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[6][3] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[6][4] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[6][5] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[6][6] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[6][7] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[7][0] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[7][1] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[7][2] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[7][3] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[7][4] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[7][5] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[7][6] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[7][7] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[8][0] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[8][1] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[8][2] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[8][3] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[8][4] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[8][5] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[8][6] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[8][7] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[9][0] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[9][1] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[9][2] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[9][3] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[9][4] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[9][5] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[9][6] ;
 wire \lut.gen_sub_units_scm.__10.sub_unit_i.mem[9][7] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.cg_we_global.clk_en ;
 wire net41;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.cg_we_global.en_i ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__0.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__1.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__10.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__11.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__12.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__13.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__14.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__15.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__16.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__17.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__18.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__19.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__2.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__20.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__21.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__22.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__23.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__24.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__25.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__26.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__27.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__28.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__29.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__3.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__30.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__31.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__4.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__5.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__6.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__7.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__8.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__9.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[0][0] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[0][1] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[0][2] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[0][3] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[0][4] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[0][5] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[0][6] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[0][7] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[10][0] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[10][1] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[10][2] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[10][3] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[10][4] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[10][5] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[10][6] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[10][7] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[11][0] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[11][1] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[11][2] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[11][3] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[11][4] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[11][5] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[11][6] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[11][7] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[12][0] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[12][1] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[12][2] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[12][3] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[12][4] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[12][5] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[12][6] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[12][7] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[13][0] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[13][1] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[13][2] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[13][3] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[13][4] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[13][5] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[13][6] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[13][7] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[14][0] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[14][1] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[14][2] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[14][3] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[14][4] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[14][5] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[14][6] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[14][7] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[15][0] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[15][1] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[15][2] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[15][3] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[15][4] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[15][5] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[15][6] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[15][7] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[16][0] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[16][1] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[16][2] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[16][3] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[16][4] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[16][5] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[16][6] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[16][7] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[17][0] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[17][1] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[17][2] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[17][3] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[17][4] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[17][5] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[17][6] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[17][7] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[18][0] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[18][1] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[18][2] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[18][3] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[18][4] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[18][5] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[18][6] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[18][7] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[19][0] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[19][1] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[19][2] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[19][3] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[19][4] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[19][5] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[19][6] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[19][7] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[1][0] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[1][1] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[1][2] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[1][3] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[1][4] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[1][5] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[1][6] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[1][7] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[20][0] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[20][1] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[20][2] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[20][3] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[20][4] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[20][5] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[20][6] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[20][7] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[21][0] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[21][1] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[21][2] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[21][3] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[21][4] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[21][5] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[21][6] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[21][7] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[22][0] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[22][1] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[22][2] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[22][3] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[22][4] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[22][5] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[22][6] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[22][7] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[23][0] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[23][1] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[23][2] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[23][3] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[23][4] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[23][5] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[23][6] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[23][7] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[24][0] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[24][1] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[24][2] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[24][3] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[24][4] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[24][5] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[24][6] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[24][7] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[25][0] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[25][1] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[25][2] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[25][3] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[25][4] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[25][5] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[25][6] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[25][7] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[26][0] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[26][1] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[26][2] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[26][3] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[26][4] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[26][5] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[26][6] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[26][7] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[27][0] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[27][1] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[27][2] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[27][3] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[27][4] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[27][5] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[27][6] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[27][7] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[28][0] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[28][1] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[28][2] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[28][3] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[28][4] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[28][5] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[28][6] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[28][7] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[29][0] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[29][1] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[29][2] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[29][3] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[29][4] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[29][5] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[29][6] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[29][7] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[2][0] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[2][1] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[2][2] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[2][3] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[2][4] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[2][5] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[2][6] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[2][7] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[30][0] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[30][1] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[30][2] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[30][3] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[30][4] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[30][5] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[30][6] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[30][7] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[31][0] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[31][1] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[31][2] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[31][3] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[31][4] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[31][5] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[31][6] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[31][7] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[3][0] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[3][1] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[3][2] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[3][3] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[3][4] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[3][5] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[3][6] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[3][7] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[4][0] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[4][1] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[4][2] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[4][3] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[4][4] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[4][5] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[4][6] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[4][7] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[5][0] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[5][1] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[5][2] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[5][3] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[5][4] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[5][5] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[5][6] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[5][7] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[6][0] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[6][1] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[6][2] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[6][3] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[6][4] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[6][5] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[6][6] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[6][7] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[7][0] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[7][1] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[7][2] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[7][3] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[7][4] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[7][5] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[7][6] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[7][7] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[8][0] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[8][1] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[8][2] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[8][3] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[8][4] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[8][5] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[8][6] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[8][7] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[9][0] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[9][1] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[9][2] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[9][3] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[9][4] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[9][5] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[9][6] ;
 wire \lut.gen_sub_units_scm.__11.sub_unit_i.mem[9][7] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.cg_we_global.clk_en ;
 wire net44;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.cg_we_global.en_i ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__0.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__1.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__10.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__11.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__12.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__13.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__14.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__15.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__16.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__17.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__18.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__19.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__2.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__20.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__21.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__22.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__23.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__24.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__25.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__26.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__27.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__28.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__29.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__3.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__30.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__31.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__4.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__5.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__6.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__7.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__8.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__9.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[0][0] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[0][1] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[0][2] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[0][3] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[0][4] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[0][5] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[0][6] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[0][7] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[10][0] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[10][1] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[10][2] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[10][3] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[10][4] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[10][5] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[10][6] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[10][7] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[11][0] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[11][1] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[11][2] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[11][3] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[11][4] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[11][5] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[11][6] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[11][7] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[12][0] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[12][1] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[12][2] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[12][3] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[12][4] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[12][5] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[12][6] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[12][7] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[13][0] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[13][1] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[13][2] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[13][3] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[13][4] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[13][5] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[13][6] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[13][7] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[14][0] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[14][1] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[14][2] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[14][3] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[14][4] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[14][5] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[14][6] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[14][7] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[15][0] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[15][1] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[15][2] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[15][3] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[15][4] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[15][5] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[15][6] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[15][7] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[16][0] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[16][1] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[16][2] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[16][3] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[16][4] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[16][5] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[16][6] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[16][7] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[17][0] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[17][1] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[17][2] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[17][3] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[17][4] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[17][5] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[17][6] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[17][7] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[18][0] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[18][1] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[18][2] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[18][3] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[18][4] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[18][5] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[18][6] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[18][7] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[19][0] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[19][1] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[19][2] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[19][3] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[19][4] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[19][5] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[19][6] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[19][7] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[1][0] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[1][1] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[1][2] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[1][3] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[1][4] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[1][5] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[1][6] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[1][7] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[20][0] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[20][1] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[20][2] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[20][3] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[20][4] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[20][5] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[20][6] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[20][7] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[21][0] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[21][1] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[21][2] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[21][3] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[21][4] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[21][5] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[21][6] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[21][7] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[22][0] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[22][1] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[22][2] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[22][3] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[22][4] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[22][5] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[22][6] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[22][7] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[23][0] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[23][1] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[23][2] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[23][3] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[23][4] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[23][5] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[23][6] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[23][7] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[24][0] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[24][1] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[24][2] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[24][3] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[24][4] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[24][5] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[24][6] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[24][7] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[25][0] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[25][1] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[25][2] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[25][3] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[25][4] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[25][5] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[25][6] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[25][7] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[26][0] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[26][1] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[26][2] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[26][3] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[26][4] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[26][5] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[26][6] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[26][7] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[27][0] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[27][1] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[27][2] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[27][3] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[27][4] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[27][5] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[27][6] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[27][7] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[28][0] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[28][1] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[28][2] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[28][3] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[28][4] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[28][5] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[28][6] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[28][7] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[29][0] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[29][1] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[29][2] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[29][3] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[29][4] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[29][5] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[29][6] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[29][7] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[2][0] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[2][1] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[2][2] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[2][3] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[2][4] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[2][5] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[2][6] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[2][7] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[30][0] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[30][1] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[30][2] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[30][3] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[30][4] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[30][5] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[30][6] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[30][7] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[31][0] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[31][1] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[31][2] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[31][3] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[31][4] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[31][5] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[31][6] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[31][7] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[3][0] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[3][1] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[3][2] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[3][3] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[3][4] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[3][5] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[3][6] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[3][7] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[4][0] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[4][1] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[4][2] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[4][3] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[4][4] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[4][5] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[4][6] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[4][7] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[5][0] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[5][1] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[5][2] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[5][3] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[5][4] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[5][5] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[5][6] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[5][7] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[6][0] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[6][1] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[6][2] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[6][3] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[6][4] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[6][5] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[6][6] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[6][7] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[7][0] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[7][1] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[7][2] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[7][3] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[7][4] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[7][5] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[7][6] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[7][7] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[8][0] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[8][1] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[8][2] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[8][3] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[8][4] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[8][5] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[8][6] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[8][7] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[9][0] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[9][1] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[9][2] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[9][3] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[9][4] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[9][5] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[9][6] ;
 wire \lut.gen_sub_units_scm.__12.sub_unit_i.mem[9][7] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.cg_we_global.clk_en ;
 wire net47;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.cg_we_global.en_i ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__0.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__1.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__10.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__11.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__12.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__13.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__14.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__15.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__16.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__17.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__18.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__19.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__2.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__20.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__21.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__22.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__23.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__24.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__25.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__26.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__27.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__28.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__29.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__3.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__30.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__31.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__4.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__5.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__6.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__7.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__8.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__9.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[0][0] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[0][1] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[0][2] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[0][3] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[0][4] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[0][5] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[0][6] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[0][7] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[10][0] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[10][1] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[10][2] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[10][3] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[10][4] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[10][5] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[10][6] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[10][7] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[11][0] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[11][1] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[11][2] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[11][3] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[11][4] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[11][5] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[11][6] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[11][7] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[12][0] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[12][1] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[12][2] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[12][3] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[12][4] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[12][5] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[12][6] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[12][7] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[13][0] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[13][1] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[13][2] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[13][3] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[13][4] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[13][5] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[13][6] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[13][7] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[14][0] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[14][1] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[14][2] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[14][3] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[14][4] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[14][5] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[14][6] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[14][7] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[15][0] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[15][1] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[15][2] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[15][3] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[15][4] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[15][5] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[15][6] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[15][7] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[16][0] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[16][1] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[16][2] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[16][3] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[16][4] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[16][5] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[16][6] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[16][7] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[17][0] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[17][1] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[17][2] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[17][3] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[17][4] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[17][5] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[17][6] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[17][7] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[18][0] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[18][1] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[18][2] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[18][3] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[18][4] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[18][5] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[18][6] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[18][7] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[19][0] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[19][1] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[19][2] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[19][3] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[19][4] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[19][5] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[19][6] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[19][7] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[1][0] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[1][1] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[1][2] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[1][3] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[1][4] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[1][5] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[1][6] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[1][7] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[20][0] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[20][1] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[20][2] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[20][3] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[20][4] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[20][5] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[20][6] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[20][7] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[21][0] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[21][1] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[21][2] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[21][3] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[21][4] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[21][5] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[21][6] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[21][7] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[22][0] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[22][1] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[22][2] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[22][3] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[22][4] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[22][5] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[22][6] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[22][7] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[23][0] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[23][1] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[23][2] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[23][3] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[23][4] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[23][5] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[23][6] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[23][7] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[24][0] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[24][1] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[24][2] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[24][3] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[24][4] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[24][5] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[24][6] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[24][7] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[25][0] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[25][1] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[25][2] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[25][3] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[25][4] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[25][5] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[25][6] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[25][7] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[26][0] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[26][1] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[26][2] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[26][3] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[26][4] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[26][5] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[26][6] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[26][7] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[27][0] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[27][1] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[27][2] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[27][3] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[27][4] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[27][5] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[27][6] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[27][7] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[28][0] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[28][1] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[28][2] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[28][3] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[28][4] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[28][5] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[28][6] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[28][7] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[29][0] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[29][1] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[29][2] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[29][3] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[29][4] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[29][5] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[29][6] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[29][7] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[2][0] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[2][1] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[2][2] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[2][3] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[2][4] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[2][5] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[2][6] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[2][7] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[30][0] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[30][1] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[30][2] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[30][3] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[30][4] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[30][5] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[30][6] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[30][7] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[31][0] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[31][1] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[31][2] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[31][3] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[31][4] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[31][5] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[31][6] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[31][7] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[3][0] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[3][1] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[3][2] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[3][3] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[3][4] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[3][5] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[3][6] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[3][7] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[4][0] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[4][1] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[4][2] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[4][3] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[4][4] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[4][5] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[4][6] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[4][7] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[5][0] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[5][1] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[5][2] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[5][3] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[5][4] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[5][5] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[5][6] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[5][7] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[6][0] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[6][1] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[6][2] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[6][3] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[6][4] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[6][5] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[6][6] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[6][7] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[7][0] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[7][1] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[7][2] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[7][3] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[7][4] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[7][5] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[7][6] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[7][7] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[8][0] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[8][1] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[8][2] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[8][3] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[8][4] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[8][5] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[8][6] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[8][7] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[9][0] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[9][1] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[9][2] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[9][3] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[9][4] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[9][5] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[9][6] ;
 wire \lut.gen_sub_units_scm.__13.sub_unit_i.mem[9][7] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.cg_we_global.clk_en ;
 wire net50;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.cg_we_global.en_i ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__0.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__1.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__10.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__11.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__12.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__13.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__14.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__15.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__16.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__17.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__18.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__19.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__2.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__20.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__21.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__22.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__23.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__24.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__25.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__26.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__27.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__28.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__29.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__3.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__30.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__31.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__4.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__5.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__6.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__7.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__8.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__9.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[0][0] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[0][1] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[0][2] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[0][3] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[0][4] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[0][5] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[0][6] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[0][7] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[10][0] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[10][1] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[10][2] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[10][3] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[10][4] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[10][5] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[10][6] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[10][7] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[11][0] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[11][1] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[11][2] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[11][3] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[11][4] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[11][5] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[11][6] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[11][7] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[12][0] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[12][1] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[12][2] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[12][3] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[12][4] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[12][5] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[12][6] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[12][7] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[13][0] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[13][1] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[13][2] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[13][3] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[13][4] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[13][5] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[13][6] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[13][7] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[14][0] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[14][1] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[14][2] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[14][3] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[14][4] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[14][5] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[14][6] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[14][7] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[15][0] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[15][1] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[15][2] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[15][3] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[15][4] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[15][5] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[15][6] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[15][7] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[16][0] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[16][1] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[16][2] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[16][3] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[16][4] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[16][5] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[16][6] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[16][7] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[17][0] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[17][1] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[17][2] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[17][3] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[17][4] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[17][5] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[17][6] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[17][7] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[18][0] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[18][1] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[18][2] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[18][3] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[18][4] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[18][5] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[18][6] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[18][7] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[19][0] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[19][1] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[19][2] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[19][3] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[19][4] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[19][5] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[19][6] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[19][7] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[1][0] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[1][1] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[1][2] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[1][3] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[1][4] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[1][5] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[1][6] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[1][7] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[20][0] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[20][1] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[20][2] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[20][3] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[20][4] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[20][5] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[20][6] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[20][7] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[21][0] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[21][1] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[21][2] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[21][3] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[21][4] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[21][5] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[21][6] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[21][7] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[22][0] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[22][1] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[22][2] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[22][3] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[22][4] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[22][5] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[22][6] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[22][7] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[23][0] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[23][1] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[23][2] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[23][3] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[23][4] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[23][5] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[23][6] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[23][7] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[24][0] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[24][1] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[24][2] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[24][3] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[24][4] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[24][5] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[24][6] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[24][7] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[25][0] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[25][1] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[25][2] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[25][3] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[25][4] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[25][5] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[25][6] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[25][7] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[26][0] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[26][1] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[26][2] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[26][3] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[26][4] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[26][5] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[26][6] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[26][7] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[27][0] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[27][1] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[27][2] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[27][3] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[27][4] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[27][5] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[27][6] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[27][7] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[28][0] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[28][1] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[28][2] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[28][3] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[28][4] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[28][5] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[28][6] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[28][7] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[29][0] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[29][1] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[29][2] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[29][3] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[29][4] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[29][5] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[29][6] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[29][7] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[2][0] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[2][1] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[2][2] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[2][3] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[2][4] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[2][5] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[2][6] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[2][7] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[30][0] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[30][1] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[30][2] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[30][3] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[30][4] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[30][5] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[30][6] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[30][7] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[31][0] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[31][1] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[31][2] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[31][3] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[31][4] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[31][5] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[31][6] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[31][7] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[3][0] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[3][1] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[3][2] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[3][3] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[3][4] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[3][5] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[3][6] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[3][7] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[4][0] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[4][1] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[4][2] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[4][3] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[4][4] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[4][5] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[4][6] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[4][7] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[5][0] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[5][1] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[5][2] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[5][3] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[5][4] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[5][5] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[5][6] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[5][7] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[6][0] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[6][1] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[6][2] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[6][3] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[6][4] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[6][5] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[6][6] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[6][7] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[7][0] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[7][1] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[7][2] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[7][3] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[7][4] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[7][5] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[7][6] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[7][7] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[8][0] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[8][1] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[8][2] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[8][3] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[8][4] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[8][5] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[8][6] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[8][7] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[9][0] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[9][1] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[9][2] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[9][3] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[9][4] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[9][5] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[9][6] ;
 wire \lut.gen_sub_units_scm.__14.sub_unit_i.mem[9][7] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.cg_we_global.clk_en ;
 wire net53;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.cg_we_global.en_i ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__0.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__1.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__10.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__11.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__12.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__13.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__14.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__15.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__16.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__17.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__18.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__19.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__2.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__20.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__21.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__22.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__23.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__24.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__25.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__26.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__27.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__28.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__29.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__3.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__30.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__31.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__4.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__5.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__6.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__7.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__8.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__9.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[0][0] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[0][1] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[0][2] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[0][3] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[0][4] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[0][5] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[0][6] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[0][7] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[10][0] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[10][1] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[10][2] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[10][3] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[10][4] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[10][5] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[10][6] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[10][7] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[11][0] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[11][1] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[11][2] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[11][3] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[11][4] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[11][5] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[11][6] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[11][7] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[12][0] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[12][1] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[12][2] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[12][3] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[12][4] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[12][5] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[12][6] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[12][7] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[13][0] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[13][1] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[13][2] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[13][3] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[13][4] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[13][5] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[13][6] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[13][7] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[14][0] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[14][1] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[14][2] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[14][3] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[14][4] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[14][5] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[14][6] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[14][7] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[15][0] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[15][1] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[15][2] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[15][3] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[15][4] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[15][5] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[15][6] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[15][7] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[16][0] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[16][1] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[16][2] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[16][3] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[16][4] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[16][5] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[16][6] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[16][7] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[17][0] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[17][1] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[17][2] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[17][3] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[17][4] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[17][5] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[17][6] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[17][7] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[18][0] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[18][1] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[18][2] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[18][3] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[18][4] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[18][5] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[18][6] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[18][7] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[19][0] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[19][1] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[19][2] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[19][3] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[19][4] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[19][5] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[19][6] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[19][7] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[1][0] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[1][1] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[1][2] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[1][3] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[1][4] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[1][5] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[1][6] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[1][7] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[20][0] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[20][1] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[20][2] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[20][3] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[20][4] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[20][5] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[20][6] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[20][7] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[21][0] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[21][1] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[21][2] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[21][3] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[21][4] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[21][5] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[21][6] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[21][7] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[22][0] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[22][1] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[22][2] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[22][3] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[22][4] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[22][5] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[22][6] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[22][7] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[23][0] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[23][1] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[23][2] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[23][3] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[23][4] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[23][5] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[23][6] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[23][7] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[24][0] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[24][1] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[24][2] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[24][3] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[24][4] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[24][5] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[24][6] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[24][7] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[25][0] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[25][1] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[25][2] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[25][3] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[25][4] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[25][5] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[25][6] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[25][7] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[26][0] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[26][1] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[26][2] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[26][3] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[26][4] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[26][5] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[26][6] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[26][7] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[27][0] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[27][1] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[27][2] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[27][3] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[27][4] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[27][5] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[27][6] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[27][7] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[28][0] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[28][1] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[28][2] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[28][3] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[28][4] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[28][5] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[28][6] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[28][7] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[29][0] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[29][1] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[29][2] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[29][3] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[29][4] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[29][5] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[29][6] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[29][7] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[2][0] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[2][1] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[2][2] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[2][3] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[2][4] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[2][5] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[2][6] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[2][7] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[30][0] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[30][1] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[30][2] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[30][3] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[30][4] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[30][5] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[30][6] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[30][7] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[31][0] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[31][1] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[31][2] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[31][3] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[31][4] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[31][5] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[31][6] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[31][7] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[3][0] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[3][1] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[3][2] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[3][3] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[3][4] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[3][5] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[3][6] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[3][7] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[4][0] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[4][1] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[4][2] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[4][3] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[4][4] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[4][5] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[4][6] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[4][7] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[5][0] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[5][1] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[5][2] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[5][3] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[5][4] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[5][5] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[5][6] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[5][7] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[6][0] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[6][1] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[6][2] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[6][3] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[6][4] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[6][5] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[6][6] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[6][7] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[7][0] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[7][1] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[7][2] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[7][3] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[7][4] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[7][5] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[7][6] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[7][7] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[8][0] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[8][1] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[8][2] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[8][3] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[8][4] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[8][5] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[8][6] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[8][7] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[9][0] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[9][1] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[9][2] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[9][3] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[9][4] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[9][5] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[9][6] ;
 wire \lut.gen_sub_units_scm.__15.sub_unit_i.mem[9][7] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.cg_we_global.clk_en ;
 wire net14;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.cg_we_global.en_i ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__0.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__1.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__10.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__11.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__12.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__13.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__14.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__15.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__16.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__17.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__18.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__19.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__2.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__20.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__21.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__22.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__23.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__24.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__25.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__26.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__27.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__28.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__29.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__3.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__30.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__31.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__4.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__5.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__6.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__7.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__8.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__9.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[0][0] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[0][1] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[0][2] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[0][3] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[0][4] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[0][5] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[0][6] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[0][7] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[10][0] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[10][1] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[10][2] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[10][3] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[10][4] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[10][5] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[10][6] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[10][7] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[11][0] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[11][1] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[11][2] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[11][3] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[11][4] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[11][5] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[11][6] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[11][7] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[12][0] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[12][1] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[12][2] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[12][3] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[12][4] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[12][5] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[12][6] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[12][7] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[13][0] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[13][1] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[13][2] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[13][3] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[13][4] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[13][5] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[13][6] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[13][7] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[14][0] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[14][1] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[14][2] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[14][3] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[14][4] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[14][5] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[14][6] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[14][7] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[15][0] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[15][1] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[15][2] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[15][3] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[15][4] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[15][5] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[15][6] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[15][7] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[16][0] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[16][1] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[16][2] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[16][3] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[16][4] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[16][5] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[16][6] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[16][7] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[17][0] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[17][1] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[17][2] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[17][3] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[17][4] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[17][5] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[17][6] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[17][7] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[18][0] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[18][1] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[18][2] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[18][3] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[18][4] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[18][5] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[18][6] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[18][7] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[19][0] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[19][1] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[19][2] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[19][3] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[19][4] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[19][5] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[19][6] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[19][7] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[1][0] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[1][1] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[1][2] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[1][3] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[1][4] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[1][5] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[1][6] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[1][7] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[20][0] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[20][1] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[20][2] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[20][3] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[20][4] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[20][5] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[20][6] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[20][7] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[21][0] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[21][1] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[21][2] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[21][3] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[21][4] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[21][5] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[21][6] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[21][7] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[22][0] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[22][1] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[22][2] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[22][3] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[22][4] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[22][5] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[22][6] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[22][7] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[23][0] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[23][1] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[23][2] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[23][3] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[23][4] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[23][5] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[23][6] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[23][7] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[24][0] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[24][1] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[24][2] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[24][3] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[24][4] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[24][5] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[24][6] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[24][7] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[25][0] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[25][1] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[25][2] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[25][3] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[25][4] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[25][5] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[25][6] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[25][7] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[26][0] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[26][1] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[26][2] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[26][3] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[26][4] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[26][5] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[26][6] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[26][7] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[27][0] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[27][1] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[27][2] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[27][3] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[27][4] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[27][5] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[27][6] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[27][7] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[28][0] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[28][1] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[28][2] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[28][3] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[28][4] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[28][5] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[28][6] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[28][7] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[29][0] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[29][1] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[29][2] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[29][3] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[29][4] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[29][5] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[29][6] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[29][7] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[2][0] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[2][1] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[2][2] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[2][3] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[2][4] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[2][5] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[2][6] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[2][7] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[30][0] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[30][1] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[30][2] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[30][3] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[30][4] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[30][5] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[30][6] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[30][7] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[31][0] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[31][1] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[31][2] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[31][3] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[31][4] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[31][5] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[31][6] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[31][7] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[3][0] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[3][1] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[3][2] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[3][3] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[3][4] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[3][5] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[3][6] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[3][7] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[4][0] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[4][1] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[4][2] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[4][3] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[4][4] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[4][5] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[4][6] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[4][7] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[5][0] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[5][1] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[5][2] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[5][3] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[5][4] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[5][5] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[5][6] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[5][7] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[6][0] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[6][1] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[6][2] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[6][3] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[6][4] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[6][5] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[6][6] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[6][7] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[7][0] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[7][1] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[7][2] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[7][3] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[7][4] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[7][5] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[7][6] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[7][7] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[8][0] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[8][1] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[8][2] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[8][3] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[8][4] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[8][5] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[8][6] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[8][7] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[9][0] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[9][1] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[9][2] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[9][3] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[9][4] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[9][5] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[9][6] ;
 wire \lut.gen_sub_units_scm.__2.sub_unit_i.mem[9][7] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.cg_we_global.clk_en ;
 wire net17;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.cg_we_global.en_i ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__0.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__1.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__10.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__11.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__12.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__13.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__14.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__15.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__16.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__17.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__18.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__19.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__2.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__20.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__21.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__22.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__23.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__24.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__25.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__26.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__27.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__28.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__29.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__3.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__30.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__31.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__4.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__5.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__6.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__7.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__8.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__9.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[0][0] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[0][1] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[0][2] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[0][3] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[0][4] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[0][5] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[0][6] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[0][7] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[10][0] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[10][1] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[10][2] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[10][3] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[10][4] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[10][5] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[10][6] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[10][7] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[11][0] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[11][1] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[11][2] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[11][3] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[11][4] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[11][5] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[11][6] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[11][7] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[12][0] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[12][1] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[12][2] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[12][3] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[12][4] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[12][5] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[12][6] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[12][7] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[13][0] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[13][1] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[13][2] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[13][3] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[13][4] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[13][5] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[13][6] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[13][7] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[14][0] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[14][1] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[14][2] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[14][3] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[14][4] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[14][5] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[14][6] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[14][7] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[15][0] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[15][1] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[15][2] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[15][3] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[15][4] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[15][5] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[15][6] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[15][7] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[16][0] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[16][1] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[16][2] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[16][3] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[16][4] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[16][5] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[16][6] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[16][7] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[17][0] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[17][1] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[17][2] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[17][3] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[17][4] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[17][5] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[17][6] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[17][7] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[18][0] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[18][1] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[18][2] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[18][3] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[18][4] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[18][5] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[18][6] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[18][7] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[19][0] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[19][1] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[19][2] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[19][3] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[19][4] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[19][5] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[19][6] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[19][7] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[1][0] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[1][1] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[1][2] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[1][3] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[1][4] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[1][5] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[1][6] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[1][7] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[20][0] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[20][1] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[20][2] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[20][3] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[20][4] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[20][5] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[20][6] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[20][7] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[21][0] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[21][1] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[21][2] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[21][3] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[21][4] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[21][5] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[21][6] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[21][7] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[22][0] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[22][1] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[22][2] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[22][3] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[22][4] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[22][5] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[22][6] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[22][7] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[23][0] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[23][1] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[23][2] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[23][3] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[23][4] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[23][5] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[23][6] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[23][7] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[24][0] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[24][1] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[24][2] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[24][3] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[24][4] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[24][5] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[24][6] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[24][7] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[25][0] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[25][1] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[25][2] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[25][3] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[25][4] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[25][5] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[25][6] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[25][7] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[26][0] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[26][1] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[26][2] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[26][3] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[26][4] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[26][5] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[26][6] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[26][7] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[27][0] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[27][1] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[27][2] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[27][3] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[27][4] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[27][5] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[27][6] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[27][7] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[28][0] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[28][1] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[28][2] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[28][3] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[28][4] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[28][5] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[28][6] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[28][7] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[29][0] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[29][1] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[29][2] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[29][3] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[29][4] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[29][5] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[29][6] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[29][7] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[2][0] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[2][1] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[2][2] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[2][3] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[2][4] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[2][5] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[2][6] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[2][7] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[30][0] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[30][1] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[30][2] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[30][3] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[30][4] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[30][5] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[30][6] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[30][7] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[31][0] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[31][1] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[31][2] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[31][3] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[31][4] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[31][5] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[31][6] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[31][7] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[3][0] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[3][1] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[3][2] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[3][3] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[3][4] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[3][5] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[3][6] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[3][7] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[4][0] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[4][1] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[4][2] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[4][3] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[4][4] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[4][5] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[4][6] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[4][7] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[5][0] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[5][1] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[5][2] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[5][3] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[5][4] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[5][5] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[5][6] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[5][7] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[6][0] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[6][1] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[6][2] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[6][3] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[6][4] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[6][5] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[6][6] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[6][7] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[7][0] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[7][1] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[7][2] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[7][3] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[7][4] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[7][5] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[7][6] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[7][7] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[8][0] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[8][1] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[8][2] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[8][3] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[8][4] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[8][5] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[8][6] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[8][7] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[9][0] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[9][1] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[9][2] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[9][3] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[9][4] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[9][5] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[9][6] ;
 wire \lut.gen_sub_units_scm.__3.sub_unit_i.mem[9][7] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.cg_we_global.clk_en ;
 wire net20;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.cg_we_global.en_i ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__0.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__1.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__10.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__11.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__12.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__13.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__14.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__15.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__16.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__17.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__18.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__19.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__2.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__20.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__21.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__22.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__23.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__24.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__25.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__26.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__27.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__28.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__29.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__3.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__30.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__31.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__4.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__5.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__6.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__7.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__8.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__9.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[0][0] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[0][1] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[0][2] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[0][3] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[0][4] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[0][5] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[0][6] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[0][7] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[10][0] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[10][1] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[10][2] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[10][3] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[10][4] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[10][5] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[10][6] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[10][7] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[11][0] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[11][1] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[11][2] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[11][3] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[11][4] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[11][5] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[11][6] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[11][7] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[12][0] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[12][1] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[12][2] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[12][3] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[12][4] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[12][5] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[12][6] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[12][7] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[13][0] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[13][1] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[13][2] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[13][3] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[13][4] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[13][5] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[13][6] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[13][7] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[14][0] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[14][1] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[14][2] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[14][3] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[14][4] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[14][5] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[14][6] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[14][7] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[15][0] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[15][1] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[15][2] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[15][3] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[15][4] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[15][5] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[15][6] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[15][7] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[16][0] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[16][1] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[16][2] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[16][3] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[16][4] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[16][5] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[16][6] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[16][7] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[17][0] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[17][1] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[17][2] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[17][3] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[17][4] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[17][5] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[17][6] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[17][7] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[18][0] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[18][1] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[18][2] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[18][3] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[18][4] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[18][5] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[18][6] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[18][7] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[19][0] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[19][1] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[19][2] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[19][3] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[19][4] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[19][5] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[19][6] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[19][7] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[1][0] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[1][1] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[1][2] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[1][3] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[1][4] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[1][5] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[1][6] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[1][7] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[20][0] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[20][1] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[20][2] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[20][3] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[20][4] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[20][5] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[20][6] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[20][7] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[21][0] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[21][1] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[21][2] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[21][3] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[21][4] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[21][5] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[21][6] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[21][7] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[22][0] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[22][1] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[22][2] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[22][3] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[22][4] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[22][5] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[22][6] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[22][7] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[23][0] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[23][1] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[23][2] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[23][3] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[23][4] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[23][5] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[23][6] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[23][7] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[24][0] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[24][1] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[24][2] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[24][3] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[24][4] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[24][5] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[24][6] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[24][7] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[25][0] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[25][1] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[25][2] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[25][3] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[25][4] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[25][5] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[25][6] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[25][7] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[26][0] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[26][1] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[26][2] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[26][3] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[26][4] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[26][5] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[26][6] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[26][7] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[27][0] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[27][1] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[27][2] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[27][3] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[27][4] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[27][5] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[27][6] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[27][7] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[28][0] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[28][1] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[28][2] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[28][3] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[28][4] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[28][5] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[28][6] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[28][7] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[29][0] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[29][1] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[29][2] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[29][3] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[29][4] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[29][5] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[29][6] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[29][7] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[2][0] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[2][1] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[2][2] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[2][3] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[2][4] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[2][5] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[2][6] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[2][7] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[30][0] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[30][1] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[30][2] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[30][3] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[30][4] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[30][5] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[30][6] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[30][7] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[31][0] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[31][1] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[31][2] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[31][3] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[31][4] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[31][5] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[31][6] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[31][7] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[3][0] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[3][1] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[3][2] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[3][3] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[3][4] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[3][5] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[3][6] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[3][7] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[4][0] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[4][1] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[4][2] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[4][3] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[4][4] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[4][5] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[4][6] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[4][7] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[5][0] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[5][1] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[5][2] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[5][3] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[5][4] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[5][5] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[5][6] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[5][7] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[6][0] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[6][1] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[6][2] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[6][3] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[6][4] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[6][5] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[6][6] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[6][7] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[7][0] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[7][1] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[7][2] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[7][3] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[7][4] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[7][5] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[7][6] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[7][7] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[8][0] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[8][1] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[8][2] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[8][3] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[8][4] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[8][5] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[8][6] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[8][7] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[9][0] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[9][1] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[9][2] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[9][3] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[9][4] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[9][5] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[9][6] ;
 wire \lut.gen_sub_units_scm.__4.sub_unit_i.mem[9][7] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.cg_we_global.clk_en ;
 wire net23;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.cg_we_global.en_i ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__0.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__1.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__10.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__11.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__12.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__13.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__14.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__15.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__16.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__17.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__18.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__19.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__2.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__20.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__21.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__22.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__23.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__24.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__25.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__26.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__27.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__28.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__29.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__3.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__30.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__31.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__4.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__5.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__6.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__7.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__8.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__9.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[0][0] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[0][1] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[0][2] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[0][3] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[0][4] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[0][5] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[0][6] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[0][7] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[10][0] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[10][1] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[10][2] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[10][3] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[10][4] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[10][5] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[10][6] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[10][7] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[11][0] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[11][1] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[11][2] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[11][3] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[11][4] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[11][5] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[11][6] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[11][7] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[12][0] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[12][1] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[12][2] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[12][3] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[12][4] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[12][5] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[12][6] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[12][7] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[13][0] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[13][1] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[13][2] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[13][3] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[13][4] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[13][5] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[13][6] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[13][7] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[14][0] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[14][1] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[14][2] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[14][3] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[14][4] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[14][5] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[14][6] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[14][7] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[15][0] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[15][1] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[15][2] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[15][3] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[15][4] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[15][5] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[15][6] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[15][7] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[16][0] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[16][1] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[16][2] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[16][3] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[16][4] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[16][5] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[16][6] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[16][7] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[17][0] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[17][1] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[17][2] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[17][3] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[17][4] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[17][5] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[17][6] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[17][7] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[18][0] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[18][1] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[18][2] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[18][3] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[18][4] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[18][5] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[18][6] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[18][7] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[19][0] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[19][1] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[19][2] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[19][3] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[19][4] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[19][5] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[19][6] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[19][7] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[1][0] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[1][1] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[1][2] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[1][3] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[1][4] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[1][5] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[1][6] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[1][7] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[20][0] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[20][1] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[20][2] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[20][3] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[20][4] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[20][5] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[20][6] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[20][7] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[21][0] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[21][1] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[21][2] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[21][3] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[21][4] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[21][5] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[21][6] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[21][7] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[22][0] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[22][1] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[22][2] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[22][3] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[22][4] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[22][5] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[22][6] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[22][7] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[23][0] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[23][1] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[23][2] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[23][3] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[23][4] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[23][5] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[23][6] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[23][7] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[24][0] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[24][1] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[24][2] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[24][3] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[24][4] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[24][5] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[24][6] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[24][7] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[25][0] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[25][1] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[25][2] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[25][3] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[25][4] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[25][5] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[25][6] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[25][7] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[26][0] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[26][1] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[26][2] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[26][3] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[26][4] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[26][5] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[26][6] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[26][7] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[27][0] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[27][1] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[27][2] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[27][3] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[27][4] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[27][5] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[27][6] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[27][7] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[28][0] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[28][1] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[28][2] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[28][3] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[28][4] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[28][5] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[28][6] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[28][7] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[29][0] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[29][1] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[29][2] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[29][3] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[29][4] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[29][5] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[29][6] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[29][7] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[2][0] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[2][1] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[2][2] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[2][3] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[2][4] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[2][5] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[2][6] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[2][7] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[30][0] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[30][1] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[30][2] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[30][3] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[30][4] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[30][5] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[30][6] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[30][7] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[31][0] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[31][1] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[31][2] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[31][3] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[31][4] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[31][5] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[31][6] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[31][7] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[3][0] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[3][1] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[3][2] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[3][3] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[3][4] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[3][5] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[3][6] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[3][7] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[4][0] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[4][1] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[4][2] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[4][3] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[4][4] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[4][5] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[4][6] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[4][7] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[5][0] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[5][1] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[5][2] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[5][3] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[5][4] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[5][5] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[5][6] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[5][7] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[6][0] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[6][1] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[6][2] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[6][3] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[6][4] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[6][5] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[6][6] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[6][7] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[7][0] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[7][1] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[7][2] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[7][3] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[7][4] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[7][5] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[7][6] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[7][7] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[8][0] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[8][1] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[8][2] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[8][3] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[8][4] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[8][5] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[8][6] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[8][7] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[9][0] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[9][1] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[9][2] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[9][3] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[9][4] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[9][5] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[9][6] ;
 wire \lut.gen_sub_units_scm.__5.sub_unit_i.mem[9][7] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.cg_we_global.clk_en ;
 wire net26;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.cg_we_global.en_i ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__0.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__1.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__10.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__11.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__12.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__13.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__14.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__15.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__16.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__17.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__18.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__19.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__2.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__20.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__21.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__22.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__23.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__24.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__25.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__26.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__27.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__28.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__29.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__3.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__30.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__31.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__4.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__5.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__6.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__7.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__8.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__9.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[0][0] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[0][1] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[0][2] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[0][3] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[0][4] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[0][5] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[0][6] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[0][7] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[10][0] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[10][1] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[10][2] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[10][3] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[10][4] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[10][5] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[10][6] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[10][7] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[11][0] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[11][1] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[11][2] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[11][3] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[11][4] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[11][5] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[11][6] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[11][7] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[12][0] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[12][1] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[12][2] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[12][3] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[12][4] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[12][5] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[12][6] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[12][7] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[13][0] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[13][1] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[13][2] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[13][3] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[13][4] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[13][5] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[13][6] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[13][7] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[14][0] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[14][1] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[14][2] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[14][3] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[14][4] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[14][5] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[14][6] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[14][7] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[15][0] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[15][1] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[15][2] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[15][3] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[15][4] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[15][5] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[15][6] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[15][7] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[16][0] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[16][1] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[16][2] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[16][3] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[16][4] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[16][5] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[16][6] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[16][7] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[17][0] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[17][1] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[17][2] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[17][3] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[17][4] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[17][5] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[17][6] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[17][7] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[18][0] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[18][1] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[18][2] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[18][3] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[18][4] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[18][5] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[18][6] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[18][7] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[19][0] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[19][1] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[19][2] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[19][3] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[19][4] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[19][5] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[19][6] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[19][7] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[1][0] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[1][1] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[1][2] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[1][3] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[1][4] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[1][5] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[1][6] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[1][7] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[20][0] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[20][1] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[20][2] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[20][3] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[20][4] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[20][5] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[20][6] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[20][7] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[21][0] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[21][1] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[21][2] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[21][3] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[21][4] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[21][5] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[21][6] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[21][7] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[22][0] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[22][1] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[22][2] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[22][3] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[22][4] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[22][5] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[22][6] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[22][7] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[23][0] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[23][1] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[23][2] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[23][3] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[23][4] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[23][5] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[23][6] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[23][7] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[24][0] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[24][1] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[24][2] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[24][3] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[24][4] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[24][5] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[24][6] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[24][7] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[25][0] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[25][1] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[25][2] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[25][3] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[25][4] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[25][5] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[25][6] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[25][7] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[26][0] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[26][1] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[26][2] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[26][3] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[26][4] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[26][5] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[26][6] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[26][7] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[27][0] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[27][1] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[27][2] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[27][3] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[27][4] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[27][5] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[27][6] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[27][7] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[28][0] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[28][1] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[28][2] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[28][3] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[28][4] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[28][5] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[28][6] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[28][7] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[29][0] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[29][1] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[29][2] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[29][3] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[29][4] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[29][5] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[29][6] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[29][7] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[2][0] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[2][1] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[2][2] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[2][3] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[2][4] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[2][5] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[2][6] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[2][7] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[30][0] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[30][1] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[30][2] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[30][3] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[30][4] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[30][5] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[30][6] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[30][7] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[31][0] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[31][1] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[31][2] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[31][3] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[31][4] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[31][5] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[31][6] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[31][7] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[3][0] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[3][1] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[3][2] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[3][3] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[3][4] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[3][5] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[3][6] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[3][7] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[4][0] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[4][1] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[4][2] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[4][3] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[4][4] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[4][5] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[4][6] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[4][7] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[5][0] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[5][1] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[5][2] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[5][3] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[5][4] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[5][5] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[5][6] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[5][7] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[6][0] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[6][1] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[6][2] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[6][3] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[6][4] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[6][5] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[6][6] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[6][7] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[7][0] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[7][1] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[7][2] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[7][3] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[7][4] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[7][5] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[7][6] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[7][7] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[8][0] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[8][1] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[8][2] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[8][3] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[8][4] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[8][5] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[8][6] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[8][7] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[9][0] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[9][1] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[9][2] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[9][3] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[9][4] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[9][5] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[9][6] ;
 wire \lut.gen_sub_units_scm.__6.sub_unit_i.mem[9][7] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.cg_we_global.clk_en ;
 wire net29;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.cg_we_global.en_i ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__0.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__1.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__10.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__11.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__12.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__13.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__14.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__15.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__16.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__17.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__18.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__19.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__2.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__20.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__21.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__22.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__23.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__24.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__25.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__26.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__27.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__28.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__29.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__3.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__30.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__31.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__4.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__5.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__6.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__7.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__8.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__9.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[0][0] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[0][1] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[0][2] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[0][3] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[0][4] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[0][5] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[0][6] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[0][7] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[10][0] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[10][1] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[10][2] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[10][3] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[10][4] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[10][5] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[10][6] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[10][7] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[11][0] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[11][1] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[11][2] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[11][3] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[11][4] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[11][5] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[11][6] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[11][7] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[12][0] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[12][1] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[12][2] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[12][3] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[12][4] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[12][5] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[12][6] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[12][7] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[13][0] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[13][1] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[13][2] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[13][3] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[13][4] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[13][5] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[13][6] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[13][7] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[14][0] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[14][1] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[14][2] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[14][3] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[14][4] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[14][5] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[14][6] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[14][7] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[15][0] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[15][1] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[15][2] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[15][3] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[15][4] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[15][5] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[15][6] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[15][7] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[16][0] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[16][1] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[16][2] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[16][3] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[16][4] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[16][5] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[16][6] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[16][7] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[17][0] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[17][1] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[17][2] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[17][3] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[17][4] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[17][5] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[17][6] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[17][7] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[18][0] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[18][1] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[18][2] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[18][3] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[18][4] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[18][5] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[18][6] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[18][7] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[19][0] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[19][1] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[19][2] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[19][3] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[19][4] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[19][5] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[19][6] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[19][7] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[1][0] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[1][1] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[1][2] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[1][3] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[1][4] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[1][5] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[1][6] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[1][7] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[20][0] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[20][1] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[20][2] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[20][3] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[20][4] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[20][5] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[20][6] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[20][7] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[21][0] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[21][1] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[21][2] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[21][3] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[21][4] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[21][5] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[21][6] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[21][7] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[22][0] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[22][1] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[22][2] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[22][3] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[22][4] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[22][5] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[22][6] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[22][7] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[23][0] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[23][1] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[23][2] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[23][3] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[23][4] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[23][5] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[23][6] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[23][7] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[24][0] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[24][1] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[24][2] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[24][3] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[24][4] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[24][5] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[24][6] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[24][7] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[25][0] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[25][1] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[25][2] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[25][3] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[25][4] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[25][5] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[25][6] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[25][7] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[26][0] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[26][1] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[26][2] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[26][3] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[26][4] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[26][5] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[26][6] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[26][7] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[27][0] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[27][1] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[27][2] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[27][3] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[27][4] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[27][5] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[27][6] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[27][7] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[28][0] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[28][1] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[28][2] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[28][3] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[28][4] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[28][5] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[28][6] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[28][7] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[29][0] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[29][1] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[29][2] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[29][3] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[29][4] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[29][5] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[29][6] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[29][7] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[2][0] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[2][1] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[2][2] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[2][3] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[2][4] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[2][5] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[2][6] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[2][7] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[30][0] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[30][1] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[30][2] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[30][3] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[30][4] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[30][5] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[30][6] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[30][7] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[31][0] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[31][1] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[31][2] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[31][3] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[31][4] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[31][5] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[31][6] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[31][7] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[3][0] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[3][1] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[3][2] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[3][3] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[3][4] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[3][5] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[3][6] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[3][7] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[4][0] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[4][1] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[4][2] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[4][3] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[4][4] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[4][5] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[4][6] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[4][7] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[5][0] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[5][1] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[5][2] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[5][3] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[5][4] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[5][5] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[5][6] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[5][7] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[6][0] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[6][1] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[6][2] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[6][3] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[6][4] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[6][5] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[6][6] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[6][7] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[7][0] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[7][1] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[7][2] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[7][3] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[7][4] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[7][5] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[7][6] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[7][7] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[8][0] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[8][1] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[8][2] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[8][3] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[8][4] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[8][5] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[8][6] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[8][7] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[9][0] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[9][1] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[9][2] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[9][3] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[9][4] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[9][5] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[9][6] ;
 wire \lut.gen_sub_units_scm.__7.sub_unit_i.mem[9][7] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.cg_we_global.clk_en ;
 wire net32;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.cg_we_global.en_i ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__0.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__1.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__10.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__11.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__12.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__13.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__14.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__15.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__16.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__17.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__18.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__19.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__2.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__20.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__21.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__22.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__23.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__24.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__25.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__26.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__27.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__28.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__29.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__3.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__30.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__31.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__4.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__5.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__6.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__7.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__8.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__9.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[0][0] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[0][1] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[0][2] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[0][3] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[0][4] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[0][5] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[0][6] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[0][7] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[10][0] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[10][1] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[10][2] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[10][3] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[10][4] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[10][5] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[10][6] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[10][7] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[11][0] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[11][1] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[11][2] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[11][3] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[11][4] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[11][5] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[11][6] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[11][7] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[12][0] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[12][1] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[12][2] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[12][3] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[12][4] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[12][5] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[12][6] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[12][7] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[13][0] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[13][1] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[13][2] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[13][3] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[13][4] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[13][5] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[13][6] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[13][7] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[14][0] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[14][1] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[14][2] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[14][3] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[14][4] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[14][5] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[14][6] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[14][7] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[15][0] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[15][1] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[15][2] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[15][3] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[15][4] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[15][5] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[15][6] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[15][7] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[16][0] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[16][1] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[16][2] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[16][3] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[16][4] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[16][5] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[16][6] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[16][7] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[17][0] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[17][1] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[17][2] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[17][3] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[17][4] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[17][5] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[17][6] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[17][7] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[18][0] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[18][1] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[18][2] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[18][3] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[18][4] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[18][5] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[18][6] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[18][7] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[19][0] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[19][1] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[19][2] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[19][3] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[19][4] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[19][5] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[19][6] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[19][7] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[1][0] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[1][1] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[1][2] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[1][3] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[1][4] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[1][5] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[1][6] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[1][7] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[20][0] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[20][1] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[20][2] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[20][3] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[20][4] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[20][5] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[20][6] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[20][7] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[21][0] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[21][1] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[21][2] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[21][3] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[21][4] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[21][5] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[21][6] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[21][7] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[22][0] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[22][1] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[22][2] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[22][3] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[22][4] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[22][5] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[22][6] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[22][7] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[23][0] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[23][1] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[23][2] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[23][3] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[23][4] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[23][5] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[23][6] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[23][7] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[24][0] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[24][1] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[24][2] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[24][3] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[24][4] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[24][5] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[24][6] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[24][7] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[25][0] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[25][1] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[25][2] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[25][3] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[25][4] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[25][5] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[25][6] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[25][7] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[26][0] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[26][1] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[26][2] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[26][3] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[26][4] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[26][5] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[26][6] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[26][7] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[27][0] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[27][1] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[27][2] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[27][3] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[27][4] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[27][5] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[27][6] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[27][7] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[28][0] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[28][1] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[28][2] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[28][3] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[28][4] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[28][5] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[28][6] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[28][7] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[29][0] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[29][1] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[29][2] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[29][3] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[29][4] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[29][5] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[29][6] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[29][7] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[2][0] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[2][1] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[2][2] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[2][3] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[2][4] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[2][5] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[2][6] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[2][7] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[30][0] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[30][1] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[30][2] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[30][3] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[30][4] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[30][5] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[30][6] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[30][7] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[31][0] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[31][1] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[31][2] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[31][3] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[31][4] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[31][5] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[31][6] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[31][7] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[3][0] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[3][1] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[3][2] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[3][3] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[3][4] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[3][5] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[3][6] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[3][7] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[4][0] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[4][1] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[4][2] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[4][3] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[4][4] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[4][5] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[4][6] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[4][7] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[5][0] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[5][1] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[5][2] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[5][3] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[5][4] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[5][5] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[5][6] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[5][7] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[6][0] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[6][1] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[6][2] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[6][3] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[6][4] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[6][5] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[6][6] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[6][7] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[7][0] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[7][1] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[7][2] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[7][3] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[7][4] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[7][5] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[7][6] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[7][7] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[8][0] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[8][1] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[8][2] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[8][3] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[8][4] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[8][5] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[8][6] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[8][7] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[9][0] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[9][1] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[9][2] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[9][3] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[9][4] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[9][5] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[9][6] ;
 wire \lut.gen_sub_units_scm.__8.sub_unit_i.mem[9][7] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.cg_we_global.clk_en ;
 wire net35;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.cg_we_global.en_i ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__0.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__1.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__10.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__11.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__12.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__13.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__14.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__15.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__16.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__17.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__18.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__19.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__2.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__20.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__21.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__22.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__23.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__24.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__25.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__26.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__27.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__28.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__29.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__3.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__30.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__31.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__4.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__5.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__6.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__7.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__8.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_en ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__9.cg_i.en_i ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[0][0] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[0][1] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[0][2] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[0][3] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[0][4] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[0][5] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[0][6] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[0][7] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[10][0] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[10][1] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[10][2] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[10][3] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[10][4] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[10][5] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[10][6] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[10][7] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[11][0] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[11][1] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[11][2] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[11][3] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[11][4] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[11][5] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[11][6] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[11][7] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[12][0] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[12][1] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[12][2] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[12][3] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[12][4] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[12][5] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[12][6] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[12][7] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[13][0] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[13][1] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[13][2] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[13][3] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[13][4] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[13][5] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[13][6] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[13][7] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[14][0] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[14][1] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[14][2] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[14][3] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[14][4] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[14][5] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[14][6] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[14][7] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[15][0] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[15][1] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[15][2] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[15][3] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[15][4] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[15][5] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[15][6] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[15][7] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[16][0] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[16][1] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[16][2] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[16][3] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[16][4] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[16][5] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[16][6] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[16][7] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[17][0] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[17][1] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[17][2] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[17][3] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[17][4] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[17][5] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[17][6] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[17][7] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[18][0] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[18][1] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[18][2] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[18][3] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[18][4] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[18][5] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[18][6] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[18][7] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[19][0] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[19][1] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[19][2] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[19][3] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[19][4] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[19][5] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[19][6] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[19][7] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[1][0] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[1][1] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[1][2] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[1][3] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[1][4] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[1][5] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[1][6] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[1][7] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[20][0] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[20][1] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[20][2] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[20][3] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[20][4] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[20][5] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[20][6] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[20][7] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[21][0] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[21][1] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[21][2] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[21][3] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[21][4] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[21][5] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[21][6] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[21][7] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[22][0] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[22][1] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[22][2] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[22][3] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[22][4] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[22][5] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[22][6] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[22][7] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[23][0] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[23][1] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[23][2] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[23][3] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[23][4] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[23][5] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[23][6] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[23][7] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[24][0] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[24][1] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[24][2] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[24][3] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[24][4] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[24][5] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[24][6] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[24][7] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[25][0] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[25][1] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[25][2] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[25][3] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[25][4] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[25][5] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[25][6] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[25][7] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[26][0] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[26][1] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[26][2] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[26][3] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[26][4] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[26][5] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[26][6] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[26][7] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[27][0] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[27][1] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[27][2] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[27][3] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[27][4] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[27][5] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[27][6] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[27][7] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[28][0] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[28][1] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[28][2] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[28][3] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[28][4] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[28][5] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[28][6] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[28][7] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[29][0] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[29][1] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[29][2] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[29][3] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[29][4] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[29][5] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[29][6] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[29][7] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[2][0] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[2][1] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[2][2] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[2][3] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[2][4] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[2][5] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[2][6] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[2][7] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[30][0] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[30][1] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[30][2] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[30][3] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[30][4] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[30][5] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[30][6] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[30][7] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[31][0] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[31][1] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[31][2] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[31][3] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[31][4] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[31][5] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[31][6] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[31][7] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[3][0] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[3][1] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[3][2] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[3][3] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[3][4] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[3][5] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[3][6] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[3][7] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[4][0] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[4][1] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[4][2] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[4][3] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[4][4] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[4][5] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[4][6] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[4][7] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[5][0] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[5][1] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[5][2] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[5][3] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[5][4] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[5][5] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[5][6] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[5][7] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[6][0] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[6][1] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[6][2] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[6][3] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[6][4] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[6][5] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[6][6] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[6][7] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[7][0] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[7][1] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[7][2] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[7][3] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[7][4] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[7][5] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[7][6] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[7][7] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[8][0] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[8][1] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[8][2] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[8][3] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[8][4] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[8][5] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[8][6] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[8][7] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[9][0] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[9][1] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[9][2] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[9][3] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[9][4] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[9][5] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[9][6] ;
 wire \lut.gen_sub_units_scm.__9.sub_unit_i.mem[9][7] ;
 wire \rdata_o_n[0] ;
 wire \rdata_o_n[1] ;
 wire \rdata_o_n[2] ;
 wire \rdata_o_n[3] ;
 wire \rdata_o_n[4] ;
 wire \rdata_o_n[5] ;
 wire \rdata_o_n[6] ;
 wire \rdata_o_n[7] ;
 wire \result_int_n[0] ;
 wire \result_int_n[10] ;
 wire \result_int_n[11] ;
 wire \result_int_n[12] ;
 wire \result_int_n[13] ;
 wire \result_int_n[14] ;
 wire \result_int_n[15] ;
 wire \result_int_n[16] ;
 wire \result_int_n[17] ;
 wire \result_int_n[18] ;
 wire \result_int_n[19] ;
 wire \result_int_n[1] ;
 wire \result_int_n[20] ;
 wire \result_int_n[21] ;
 wire \result_int_n[22] ;
 wire \result_int_n[23] ;
 wire \result_int_n[24] ;
 wire \result_int_n[25] ;
 wire \result_int_n[26] ;
 wire \result_int_n[27] ;
 wire \result_int_n[28] ;
 wire \result_int_n[29] ;
 wire \result_int_n[2] ;
 wire \result_int_n[30] ;
 wire \result_int_n[31] ;
 wire \result_int_n[3] ;
 wire \result_int_n[4] ;
 wire \result_int_n[5] ;
 wire \result_int_n[6] ;
 wire \result_int_n[7] ;
 wire \result_int_n[8] ;
 wire \result_int_n[9] ;
 wire \clknet_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ;
 wire clknet_0__00540_;
 wire clknet_3_0__leaf__00540_;
 wire clknet_3_1__leaf__00540_;
 wire clknet_3_2__leaf__00540_;
 wire clknet_3_3__leaf__00540_;
 wire clknet_3_4__leaf__00540_;
 wire clknet_3_5__leaf__00540_;
 wire clknet_3_6__leaf__00540_;
 wire clknet_3_7__leaf__00540_;
 wire clknet_level_0_1_1321__00540_;
 wire clknet_level_1_1_1322__00540_;
 wire clknet_level_2_1_1323__00540_;
 wire clknet_level_0_1_2324__00540_;
 wire clknet_level_1_1_2325__00540_;
 wire clknet_level_2_1_2326__00540_;
 wire clknet_level_0_1_3327__00540_;
 wire clknet_level_1_1_3328__00540_;
 wire clknet_level_2_1_3329__00540_;
 wire clknet_level_0_1_4330__00540_;
 wire clknet_level_1_1_4331__00540_;
 wire clknet_level_2_1_4332__00540_;
 wire clknet_level_0_1_5333__00540_;
 wire clknet_level_1_1_5334__00540_;
 wire clknet_level_2_1_5335__00540_;
 wire clknet_level_0_1_6336__00540_;
 wire clknet_level_1_1_6337__00540_;
 wire clknet_level_2_1_6338__00540_;
 wire clknet_level_0_1_7339__00540_;
 wire clknet_level_1_1_7340__00540_;
 wire clknet_level_2_1_7341__00540_;
 wire clknet_level_0_1_8342__00540_;
 wire clknet_level_1_1_8343__00540_;
 wire clknet_level_2_1_8344__00540_;
 wire \clknet_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ;
 wire clknet_0__00543_;
 wire clknet_3_0__leaf__00543_;
 wire clknet_3_1__leaf__00543_;
 wire clknet_3_2__leaf__00543_;
 wire clknet_3_3__leaf__00543_;
 wire clknet_3_4__leaf__00543_;
 wire clknet_3_5__leaf__00543_;
 wire clknet_3_6__leaf__00543_;
 wire clknet_3_7__leaf__00543_;
 wire clknet_level_0_1_1141__00543_;
 wire clknet_level_1_1_1142__00543_;
 wire clknet_level_2_1_1143__00543_;
 wire clknet_level_0_1_2144__00543_;
 wire clknet_level_1_1_2145__00543_;
 wire clknet_level_2_1_2146__00543_;
 wire clknet_level_0_1_3147__00543_;
 wire clknet_level_1_1_3148__00543_;
 wire clknet_level_2_1_3149__00543_;
 wire clknet_level_0_1_4150__00543_;
 wire clknet_level_1_1_4151__00543_;
 wire clknet_level_2_1_4152__00543_;
 wire clknet_level_0_1_5153__00543_;
 wire clknet_level_1_1_5154__00543_;
 wire clknet_level_2_1_5155__00543_;
 wire clknet_level_0_1_6156__00543_;
 wire clknet_level_1_1_6157__00543_;
 wire clknet_level_2_1_6158__00543_;
 wire clknet_level_0_1_7159__00543_;
 wire clknet_level_1_1_7160__00543_;
 wire clknet_level_2_1_7161__00543_;
 wire clknet_level_0_1_8162__00543_;
 wire clknet_level_1_1_8163__00543_;
 wire clknet_level_2_1_8164__00543_;
 wire \clknet_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ;
 wire clknet_0__00546_;
 wire clknet_3_0__leaf__00546_;
 wire clknet_3_1__leaf__00546_;
 wire clknet_3_2__leaf__00546_;
 wire clknet_3_3__leaf__00546_;
 wire clknet_3_4__leaf__00546_;
 wire clknet_3_5__leaf__00546_;
 wire clknet_3_6__leaf__00546_;
 wire clknet_3_7__leaf__00546_;
 wire clknet_level_0_1_1345__00546_;
 wire clknet_level_1_1_1346__00546_;
 wire clknet_level_2_1_1347__00546_;
 wire clknet_level_0_1_2348__00546_;
 wire clknet_level_1_1_2349__00546_;
 wire clknet_level_2_1_2350__00546_;
 wire clknet_level_0_1_3351__00546_;
 wire clknet_level_1_1_3352__00546_;
 wire clknet_level_2_1_3353__00546_;
 wire clknet_level_0_1_4354__00546_;
 wire clknet_level_1_1_4355__00546_;
 wire clknet_level_2_1_4356__00546_;
 wire clknet_level_0_1_5357__00546_;
 wire clknet_level_1_1_5358__00546_;
 wire clknet_level_2_1_5359__00546_;
 wire clknet_level_0_1_6360__00546_;
 wire clknet_level_1_1_6361__00546_;
 wire clknet_level_2_1_6362__00546_;
 wire clknet_level_0_1_7363__00546_;
 wire clknet_level_1_1_7364__00546_;
 wire clknet_level_2_1_7365__00546_;
 wire clknet_level_0_1_8366__00546_;
 wire clknet_level_1_1_8367__00546_;
 wire clknet_level_2_1_8368__00546_;
 wire \clknet_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ;
 wire clknet_0__00549_;
 wire clknet_3_0__leaf__00549_;
 wire clknet_3_1__leaf__00549_;
 wire clknet_3_2__leaf__00549_;
 wire clknet_3_3__leaf__00549_;
 wire clknet_3_4__leaf__00549_;
 wire clknet_3_5__leaf__00549_;
 wire clknet_3_6__leaf__00549_;
 wire clknet_3_7__leaf__00549_;
 wire clknet_level_0_1_115__00549_;
 wire clknet_level_1_1_116__00549_;
 wire clknet_level_2_1_117__00549_;
 wire clknet_level_0_1_218__00549_;
 wire clknet_level_1_1_219__00549_;
 wire clknet_level_2_1_220__00549_;
 wire clknet_level_0_1_321__00549_;
 wire clknet_level_1_1_322__00549_;
 wire clknet_level_2_1_323__00549_;
 wire clknet_level_0_1_424__00549_;
 wire clknet_level_1_1_425__00549_;
 wire clknet_level_2_1_426__00549_;
 wire clknet_level_0_1_527__00549_;
 wire clknet_level_1_1_528__00549_;
 wire clknet_level_2_1_529__00549_;
 wire clknet_level_0_1_630__00549_;
 wire clknet_level_1_1_631__00549_;
 wire clknet_level_2_1_632__00549_;
 wire clknet_level_0_1_733__00549_;
 wire clknet_level_1_1_734__00549_;
 wire clknet_level_2_1_735__00549_;
 wire clknet_level_0_1_836__00549_;
 wire clknet_level_1_1_837__00549_;
 wire clknet_level_2_1_838__00549_;
 wire \clknet_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ;
 wire clknet_0__00552_;
 wire clknet_3_0__leaf__00552_;
 wire clknet_3_1__leaf__00552_;
 wire clknet_3_2__leaf__00552_;
 wire clknet_3_3__leaf__00552_;
 wire clknet_3_4__leaf__00552_;
 wire clknet_3_5__leaf__00552_;
 wire clknet_3_6__leaf__00552_;
 wire clknet_3_7__leaf__00552_;
 wire clknet_level_0_1_1165__00552_;
 wire clknet_level_1_1_1166__00552_;
 wire clknet_level_2_1_1167__00552_;
 wire clknet_level_0_1_2168__00552_;
 wire clknet_level_1_1_2169__00552_;
 wire clknet_level_2_1_2170__00552_;
 wire clknet_level_0_1_3171__00552_;
 wire clknet_level_1_1_3172__00552_;
 wire clknet_level_2_1_3173__00552_;
 wire clknet_level_0_1_4174__00552_;
 wire clknet_level_1_1_4175__00552_;
 wire clknet_level_2_1_4176__00552_;
 wire clknet_level_0_1_5177__00552_;
 wire clknet_level_1_1_5178__00552_;
 wire clknet_level_2_1_5179__00552_;
 wire clknet_level_0_1_6180__00552_;
 wire clknet_level_1_1_6181__00552_;
 wire clknet_level_2_1_6182__00552_;
 wire clknet_level_0_1_7183__00552_;
 wire clknet_level_1_1_7184__00552_;
 wire clknet_level_2_1_7185__00552_;
 wire clknet_level_0_1_8186__00552_;
 wire clknet_level_1_1_8187__00552_;
 wire clknet_level_2_1_8188__00552_;
 wire \clknet_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ;
 wire clknet_0__00555_;
 wire clknet_3_0__leaf__00555_;
 wire clknet_3_1__leaf__00555_;
 wire clknet_3_2__leaf__00555_;
 wire clknet_3_3__leaf__00555_;
 wire clknet_3_4__leaf__00555_;
 wire clknet_3_5__leaf__00555_;
 wire clknet_3_6__leaf__00555_;
 wire clknet_3_7__leaf__00555_;
 wire clknet_level_0_1_139__00555_;
 wire clknet_level_1_1_140__00555_;
 wire clknet_level_2_1_141__00555_;
 wire clknet_level_0_1_242__00555_;
 wire clknet_level_1_1_243__00555_;
 wire clknet_level_2_1_244__00555_;
 wire clknet_level_0_1_345__00555_;
 wire clknet_level_1_1_346__00555_;
 wire clknet_level_2_1_347__00555_;
 wire clknet_level_0_1_448__00555_;
 wire clknet_level_1_1_449__00555_;
 wire clknet_level_2_1_450__00555_;
 wire clknet_level_0_1_551__00555_;
 wire clknet_level_1_1_552__00555_;
 wire clknet_level_2_1_553__00555_;
 wire clknet_level_0_1_654__00555_;
 wire clknet_level_1_1_655__00555_;
 wire clknet_level_2_1_656__00555_;
 wire clknet_level_0_1_757__00555_;
 wire clknet_level_1_1_758__00555_;
 wire clknet_level_2_1_759__00555_;
 wire clknet_level_0_1_860__00555_;
 wire clknet_level_1_1_861__00555_;
 wire clknet_level_2_1_862__00555_;
 wire \clknet_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ;
 wire clknet_0__00558_;
 wire clknet_3_0__leaf__00558_;
 wire clknet_3_1__leaf__00558_;
 wire clknet_3_2__leaf__00558_;
 wire clknet_3_3__leaf__00558_;
 wire clknet_3_4__leaf__00558_;
 wire clknet_3_5__leaf__00558_;
 wire clknet_3_6__leaf__00558_;
 wire clknet_3_7__leaf__00558_;
 wire clknet_level_0_1_163__00558_;
 wire clknet_level_1_1_164__00558_;
 wire clknet_level_2_1_165__00558_;
 wire clknet_level_0_1_266__00558_;
 wire clknet_level_1_1_267__00558_;
 wire clknet_level_2_1_268__00558_;
 wire clknet_level_0_1_369__00558_;
 wire clknet_level_1_1_370__00558_;
 wire clknet_level_2_1_371__00558_;
 wire clknet_level_0_1_472__00558_;
 wire clknet_level_1_1_473__00558_;
 wire clknet_level_2_1_474__00558_;
 wire clknet_level_0_1_575__00558_;
 wire clknet_level_1_1_576__00558_;
 wire clknet_level_2_1_577__00558_;
 wire clknet_level_0_1_678__00558_;
 wire clknet_level_1_1_679__00558_;
 wire clknet_level_2_1_680__00558_;
 wire clknet_level_0_1_781__00558_;
 wire clknet_level_1_1_782__00558_;
 wire clknet_level_2_1_783__00558_;
 wire clknet_level_0_1_884__00558_;
 wire clknet_level_1_1_885__00558_;
 wire clknet_level_2_1_886__00558_;
 wire \clknet_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ;
 wire clknet_0__00561_;
 wire clknet_3_0__leaf__00561_;
 wire clknet_3_1__leaf__00561_;
 wire clknet_3_2__leaf__00561_;
 wire clknet_3_3__leaf__00561_;
 wire clknet_3_4__leaf__00561_;
 wire clknet_3_5__leaf__00561_;
 wire clknet_3_6__leaf__00561_;
 wire clknet_3_7__leaf__00561_;
 wire clknet_level_0_1_187__00561_;
 wire clknet_level_1_1_188__00561_;
 wire clknet_level_2_1_189__00561_;
 wire clknet_level_0_1_290__00561_;
 wire clknet_level_1_1_291__00561_;
 wire clknet_level_2_1_292__00561_;
 wire clknet_level_0_1_393__00561_;
 wire clknet_level_1_1_394__00561_;
 wire clknet_level_2_1_395__00561_;
 wire clknet_level_0_1_496__00561_;
 wire clknet_level_1_1_497__00561_;
 wire clknet_level_2_1_498__00561_;
 wire clknet_level_0_1_599__00561_;
 wire clknet_level_1_1_5100__00561_;
 wire clknet_level_2_1_5101__00561_;
 wire clknet_level_0_1_6102__00561_;
 wire clknet_level_1_1_6103__00561_;
 wire clknet_level_2_1_6104__00561_;
 wire clknet_level_0_1_7105__00561_;
 wire clknet_level_1_1_7106__00561_;
 wire clknet_level_2_1_7107__00561_;
 wire clknet_level_0_1_8108__00561_;
 wire clknet_level_1_1_8109__00561_;
 wire clknet_level_2_1_8110__00561_;
 wire \clknet_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ;
 wire clknet_0__00564_;
 wire clknet_3_0__leaf__00564_;
 wire clknet_3_1__leaf__00564_;
 wire clknet_3_2__leaf__00564_;
 wire clknet_3_3__leaf__00564_;
 wire clknet_3_4__leaf__00564_;
 wire clknet_3_5__leaf__00564_;
 wire clknet_3_6__leaf__00564_;
 wire clknet_3_7__leaf__00564_;
 wire clknet_level_0_1_1243__00564_;
 wire clknet_level_1_1_1244__00564_;
 wire clknet_level_2_1_1245__00564_;
 wire clknet_level_0_1_2246__00564_;
 wire clknet_level_1_1_2247__00564_;
 wire clknet_level_2_1_2248__00564_;
 wire clknet_level_0_1_3249__00564_;
 wire clknet_level_1_1_3250__00564_;
 wire clknet_level_2_1_3251__00564_;
 wire clknet_level_0_1_4252__00564_;
 wire clknet_level_1_1_4253__00564_;
 wire clknet_level_2_1_4254__00564_;
 wire clknet_level_0_1_5255__00564_;
 wire clknet_level_1_1_5256__00564_;
 wire clknet_level_2_1_5257__00564_;
 wire clknet_level_0_1_6258__00564_;
 wire clknet_level_1_1_6259__00564_;
 wire clknet_level_2_1_6260__00564_;
 wire clknet_level_0_1_7261__00564_;
 wire clknet_level_1_1_7262__00564_;
 wire clknet_level_2_1_7263__00564_;
 wire clknet_level_0_1_8264__00564_;
 wire clknet_level_1_1_8265__00564_;
 wire clknet_level_2_1_8266__00564_;
 wire \clknet_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ;
 wire clknet_0__00567_;
 wire clknet_3_0__leaf__00567_;
 wire clknet_3_1__leaf__00567_;
 wire clknet_3_2__leaf__00567_;
 wire clknet_3_3__leaf__00567_;
 wire clknet_3_4__leaf__00567_;
 wire clknet_3_5__leaf__00567_;
 wire clknet_3_6__leaf__00567_;
 wire clknet_3_7__leaf__00567_;
 wire clknet_level_0_1_1189__00567_;
 wire clknet_level_1_1_1190__00567_;
 wire clknet_level_2_1_1191__00567_;
 wire clknet_level_0_1_2192__00567_;
 wire clknet_level_1_1_2193__00567_;
 wire clknet_level_2_1_2194__00567_;
 wire clknet_level_0_1_3195__00567_;
 wire clknet_level_1_1_3196__00567_;
 wire clknet_level_2_1_3197__00567_;
 wire clknet_level_0_1_4198__00567_;
 wire clknet_level_1_1_4199__00567_;
 wire clknet_level_2_1_4200__00567_;
 wire clknet_level_0_1_5201__00567_;
 wire clknet_level_1_1_5202__00567_;
 wire clknet_level_2_1_5203__00567_;
 wire clknet_level_0_1_6204__00567_;
 wire clknet_level_1_1_6205__00567_;
 wire clknet_level_2_1_6206__00567_;
 wire clknet_level_0_1_7207__00567_;
 wire clknet_level_1_1_7208__00567_;
 wire clknet_level_2_1_7209__00567_;
 wire clknet_level_0_1_8210__00567_;
 wire clknet_level_1_1_8211__00567_;
 wire clknet_level_2_1_8212__00567_;
 wire \clknet_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ;
 wire clknet_0__00570_;
 wire clknet_3_0__leaf__00570_;
 wire clknet_3_1__leaf__00570_;
 wire clknet_3_2__leaf__00570_;
 wire clknet_3_3__leaf__00570_;
 wire clknet_3_4__leaf__00570_;
 wire clknet_3_5__leaf__00570_;
 wire clknet_3_6__leaf__00570_;
 wire clknet_3_7__leaf__00570_;
 wire clknet_level_0_1_1267__00570_;
 wire clknet_level_1_1_1268__00570_;
 wire clknet_level_2_1_1269__00570_;
 wire clknet_level_0_1_2270__00570_;
 wire clknet_level_1_1_2271__00570_;
 wire clknet_level_2_1_2272__00570_;
 wire clknet_level_0_1_3273__00570_;
 wire clknet_level_1_1_3274__00570_;
 wire clknet_level_2_1_3275__00570_;
 wire clknet_level_0_1_4276__00570_;
 wire clknet_level_1_1_4277__00570_;
 wire clknet_level_2_1_4278__00570_;
 wire clknet_level_0_1_5279__00570_;
 wire clknet_level_1_1_5280__00570_;
 wire clknet_level_2_1_5281__00570_;
 wire clknet_level_0_1_6282__00570_;
 wire clknet_level_1_1_6283__00570_;
 wire clknet_level_2_1_6284__00570_;
 wire clknet_level_0_1_7285__00570_;
 wire clknet_level_1_1_7286__00570_;
 wire clknet_level_2_1_7287__00570_;
 wire clknet_level_0_1_8288__00570_;
 wire clknet_level_1_1_8289__00570_;
 wire clknet_level_2_1_8290__00570_;
 wire \clknet_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ;
 wire clknet_0__00573_;
 wire clknet_3_0__leaf__00573_;
 wire clknet_3_1__leaf__00573_;
 wire clknet_3_2__leaf__00573_;
 wire clknet_3_3__leaf__00573_;
 wire clknet_3_4__leaf__00573_;
 wire clknet_3_5__leaf__00573_;
 wire clknet_3_6__leaf__00573_;
 wire clknet_3_7__leaf__00573_;
 wire clknet_level_0_1_1291__00573_;
 wire clknet_level_1_1_1292__00573_;
 wire clknet_level_2_1_1293__00573_;
 wire clknet_level_0_1_2294__00573_;
 wire clknet_level_1_1_2295__00573_;
 wire clknet_level_2_1_2296__00573_;
 wire clknet_level_0_1_3297__00573_;
 wire clknet_level_1_1_3298__00573_;
 wire clknet_level_2_1_3299__00573_;
 wire clknet_level_0_1_4300__00573_;
 wire clknet_level_1_1_4301__00573_;
 wire clknet_level_2_1_4302__00573_;
 wire clknet_level_0_1_5303__00573_;
 wire clknet_level_1_1_5304__00573_;
 wire clknet_level_2_1_5305__00573_;
 wire clknet_level_0_1_6306__00573_;
 wire clknet_level_1_1_6307__00573_;
 wire clknet_level_2_1_6308__00573_;
 wire clknet_level_0_1_7309__00573_;
 wire clknet_level_1_1_7310__00573_;
 wire clknet_level_2_1_7311__00573_;
 wire clknet_level_0_1_8312__00573_;
 wire clknet_level_1_1_8313__00573_;
 wire clknet_level_2_1_8314__00573_;
 wire \clknet_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ;
 wire clknet_0__00576_;
 wire clknet_3_0__leaf__00576_;
 wire clknet_3_1__leaf__00576_;
 wire clknet_3_2__leaf__00576_;
 wire clknet_3_3__leaf__00576_;
 wire clknet_3_4__leaf__00576_;
 wire clknet_3_5__leaf__00576_;
 wire clknet_3_6__leaf__00576_;
 wire clknet_3_7__leaf__00576_;
 wire clknet_level_0_1_1369__00576_;
 wire clknet_level_1_1_1370__00576_;
 wire clknet_level_2_1_1371__00576_;
 wire clknet_level_0_1_2372__00576_;
 wire clknet_level_1_1_2373__00576_;
 wire clknet_level_2_1_2374__00576_;
 wire clknet_level_0_1_3375__00576_;
 wire clknet_level_1_1_3376__00576_;
 wire clknet_level_2_1_3377__00576_;
 wire clknet_level_0_1_4378__00576_;
 wire clknet_level_1_1_4379__00576_;
 wire clknet_level_2_1_4380__00576_;
 wire clknet_level_0_1_5381__00576_;
 wire clknet_level_1_1_5382__00576_;
 wire clknet_level_2_1_5383__00576_;
 wire clknet_level_0_1_6384__00576_;
 wire clknet_level_1_1_6385__00576_;
 wire clknet_level_2_1_6386__00576_;
 wire clknet_level_0_1_7387__00576_;
 wire clknet_level_1_1_7388__00576_;
 wire clknet_level_2_1_7389__00576_;
 wire clknet_level_0_1_8390__00576_;
 wire clknet_level_1_1_8391__00576_;
 wire clknet_level_2_1_8392__00576_;
 wire \clknet_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ;
 wire clknet_0__00579_;
 wire clknet_3_0__leaf__00579_;
 wire clknet_3_1__leaf__00579_;
 wire clknet_3_2__leaf__00579_;
 wire clknet_3_3__leaf__00579_;
 wire clknet_3_4__leaf__00579_;
 wire clknet_3_5__leaf__00579_;
 wire clknet_3_6__leaf__00579_;
 wire clknet_3_7__leaf__00579_;
 wire clknet_level_0_1_1393__00579_;
 wire clknet_level_1_1_1394__00579_;
 wire clknet_level_2_1_1395__00579_;
 wire clknet_level_0_1_2396__00579_;
 wire clknet_level_1_1_2397__00579_;
 wire clknet_level_2_1_2398__00579_;
 wire clknet_level_0_1_3399__00579_;
 wire clknet_level_1_1_3400__00579_;
 wire clknet_level_2_1_3401__00579_;
 wire clknet_level_0_1_4402__00579_;
 wire clknet_level_1_1_4403__00579_;
 wire clknet_level_2_1_4404__00579_;
 wire clknet_level_0_1_5405__00579_;
 wire clknet_level_1_1_5406__00579_;
 wire clknet_level_2_1_5407__00579_;
 wire clknet_level_0_1_6408__00579_;
 wire clknet_level_1_1_6409__00579_;
 wire clknet_level_2_1_6410__00579_;
 wire clknet_level_0_1_7411__00579_;
 wire clknet_level_1_1_7412__00579_;
 wire clknet_level_2_1_7413__00579_;
 wire clknet_level_0_1_8414__00579_;
 wire clknet_level_1_1_8415__00579_;
 wire clknet_level_2_1_8416__00579_;
 wire \clknet_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ;
 wire \clknet_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ;
 wire \clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ;
 wire \clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ;

 BUF_X4 max_cap231 (.A(_00993_),
    .Z(net231));
 BUF_X4 max_cap230 (.A(_00993_),
    .Z(net230));
 BUF_X8 max_cap229 (.A(net230),
    .Z(net229));
 BUF_X8 max_cap228 (.A(_00996_),
    .Z(net228));
 AND3_X4 _04314_ (.A1(net20),
    .A2(net19),
    .A3(net29),
    .ZN(_00655_));
 NAND3_X4 _04315_ (.A1(net18),
    .A2(net17),
    .A3(_00655_),
    .ZN(_00656_));
 BUF_X8 max_cap227 (.A(_00996_),
    .Z(net227));
 INV_X1 _04317_ (.A(_00656_),
    .ZN(\lut.gen_sub_units_scm.__15.sub_unit_i.cg_we_global.en_i ));
 BUF_X8 wire226 (.A(_00996_),
    .Z(net226));
 BUF_X16 max_cap225 (.A(net226),
    .Z(net225));
 NOR2_X1 _04320_ (.A1(net16),
    .A2(net12),
    .ZN(_00660_));
 BUF_X8 max_cap224 (.A(net225),
    .Z(net224));
 BUF_X8 max_cap223 (.A(net225),
    .Z(net223));
 BUF_X8 max_cap222 (.A(net226),
    .Z(net222));
 NOR3_X4 _04324_ (.A1(net13),
    .A2(net14),
    .A3(net15),
    .ZN(_00664_));
 NAND2_X4 _04325_ (.A1(_00660_),
    .A2(_00664_),
    .ZN(_00665_));
 NOR2_X1 _04326_ (.A1(_00656_),
    .A2(_00665_),
    .ZN(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__0.cg_i.en_i ));
 INV_X2 _04327_ (.A(net12),
    .ZN(_00666_));
 NOR2_X1 _04328_ (.A1(net16),
    .A2(_00666_),
    .ZN(_00667_));
 NAND2_X4 _04329_ (.A1(_00664_),
    .A2(_00667_),
    .ZN(_00668_));
 NOR2_X1 _04330_ (.A1(_00656_),
    .A2(_00668_),
    .ZN(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__1.cg_i.en_i ));
 NOR2_X4 _04331_ (.A1(net14),
    .A2(net15),
    .ZN(_00669_));
 AND2_X2 _04332_ (.A1(net13),
    .A2(_00660_),
    .ZN(_00670_));
 NAND2_X4 _04333_ (.A1(_00669_),
    .A2(_00670_),
    .ZN(_00671_));
 NOR2_X1 _04334_ (.A1(_00656_),
    .A2(_00671_),
    .ZN(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__2.cg_i.en_i ));
 AND2_X2 _04335_ (.A1(net13),
    .A2(_00667_),
    .ZN(_00672_));
 NAND2_X4 _04336_ (.A1(_00669_),
    .A2(_00672_),
    .ZN(_00673_));
 NOR2_X1 _04337_ (.A1(_00656_),
    .A2(_00673_),
    .ZN(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__3.cg_i.en_i ));
 INV_X2 _04338_ (.A(net14),
    .ZN(_00674_));
 NOR2_X4 _04339_ (.A1(_00674_),
    .A2(net15),
    .ZN(_00675_));
 BUF_X8 max_cap221 (.A(_00999_),
    .Z(net221));
 NOR3_X4 _04341_ (.A1(net16),
    .A2(net12),
    .A3(net13),
    .ZN(_00677_));
 NAND2_X4 _04342_ (.A1(_00675_),
    .A2(_00677_),
    .ZN(_00678_));
 NOR2_X1 _04343_ (.A1(_00656_),
    .A2(_00678_),
    .ZN(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__4.cg_i.en_i ));
 NOR3_X4 _04344_ (.A1(net16),
    .A2(_00666_),
    .A3(net13),
    .ZN(_00679_));
 NAND2_X4 _04345_ (.A1(_00675_),
    .A2(_00679_),
    .ZN(_00680_));
 NOR2_X1 _04346_ (.A1(_00656_),
    .A2(_00680_),
    .ZN(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__5.cg_i.en_i ));
 NAND2_X4 _04347_ (.A1(_00670_),
    .A2(_00675_),
    .ZN(_00681_));
 NOR2_X1 _04348_ (.A1(_00656_),
    .A2(_00681_),
    .ZN(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__6.cg_i.en_i ));
 NAND2_X4 _04349_ (.A1(_00672_),
    .A2(_00675_),
    .ZN(_00682_));
 NOR2_X1 _04350_ (.A1(_00656_),
    .A2(_00682_),
    .ZN(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__7.cg_i.en_i ));
 INV_X2 _04351_ (.A(net15),
    .ZN(_00683_));
 NOR2_X4 _04352_ (.A1(net14),
    .A2(_00683_),
    .ZN(_00684_));
 BUF_X8 wire220 (.A(net221),
    .Z(net220));
 NAND2_X4 _04354_ (.A1(_00677_),
    .A2(_00684_),
    .ZN(_00686_));
 NOR2_X1 _04355_ (.A1(_00656_),
    .A2(_00686_),
    .ZN(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__8.cg_i.en_i ));
 BUF_X8 max_cap219 (.A(net220),
    .Z(net219));
 NAND2_X4 _04357_ (.A1(_00679_),
    .A2(_00684_),
    .ZN(_00688_));
 NOR2_X1 _04358_ (.A1(_00656_),
    .A2(_00688_),
    .ZN(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__9.cg_i.en_i ));
 NAND2_X4 _04359_ (.A1(_00670_),
    .A2(_00684_),
    .ZN(_00689_));
 NOR2_X1 _04360_ (.A1(_00656_),
    .A2(_00689_),
    .ZN(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__10.cg_i.en_i ));
 NAND2_X4 _04361_ (.A1(_00672_),
    .A2(_00684_),
    .ZN(_00690_));
 NOR2_X1 _04362_ (.A1(_00656_),
    .A2(_00690_),
    .ZN(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__11.cg_i.en_i ));
 NOR2_X4 _04363_ (.A1(_00674_),
    .A2(_00683_),
    .ZN(_00691_));
 BUF_X8 max_cap218 (.A(net221),
    .Z(net218));
 NAND2_X4 _04365_ (.A1(_00677_),
    .A2(_00691_),
    .ZN(_00693_));
 NOR2_X1 _04366_ (.A1(_00656_),
    .A2(_00693_),
    .ZN(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__12.cg_i.en_i ));
 NAND2_X4 _04367_ (.A1(_00679_),
    .A2(_00691_),
    .ZN(_00694_));
 NOR2_X1 _04368_ (.A1(_00656_),
    .A2(_00694_),
    .ZN(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__13.cg_i.en_i ));
 NAND2_X4 _04369_ (.A1(_00670_),
    .A2(_00691_),
    .ZN(_00695_));
 NOR2_X1 _04370_ (.A1(_00656_),
    .A2(_00695_),
    .ZN(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__14.cg_i.en_i ));
 NAND2_X4 _04371_ (.A1(_00672_),
    .A2(_00691_),
    .ZN(_00696_));
 NOR2_X1 _04372_ (.A1(_00656_),
    .A2(_00696_),
    .ZN(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__15.cg_i.en_i ));
 INV_X2 _04373_ (.A(net16),
    .ZN(_00697_));
 NOR2_X1 _04374_ (.A1(_00697_),
    .A2(net12),
    .ZN(_00698_));
 NAND2_X4 _04375_ (.A1(_00664_),
    .A2(_00698_),
    .ZN(_00699_));
 NOR2_X1 _04376_ (.A1(_00656_),
    .A2(_00699_),
    .ZN(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__16.cg_i.en_i ));
 NAND3_X4 _04377_ (.A1(net16),
    .A2(net12),
    .A3(_00664_),
    .ZN(_00700_));
 NOR2_X1 _04378_ (.A1(_00656_),
    .A2(_00700_),
    .ZN(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__17.cg_i.en_i ));
 AND2_X2 _04379_ (.A1(net13),
    .A2(_00698_),
    .ZN(_00701_));
 BUF_X8 max_cap217 (.A(net218),
    .Z(net217));
 NAND2_X4 _04381_ (.A1(_00669_),
    .A2(_00701_),
    .ZN(_00703_));
 NOR2_X1 _04382_ (.A1(_00656_),
    .A2(_00703_),
    .ZN(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__18.cg_i.en_i ));
 BUF_X4 max_cap216 (.A(_01002_),
    .Z(net216));
 AND3_X4 _04384_ (.A1(net16),
    .A2(net12),
    .A3(net13),
    .ZN(_00705_));
 BUF_X8 max_cap215 (.A(net216),
    .Z(net215));
 NAND2_X4 _04386_ (.A1(_00669_),
    .A2(_00705_),
    .ZN(_00707_));
 NOR2_X1 _04387_ (.A1(_00656_),
    .A2(_00707_),
    .ZN(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__19.cg_i.en_i ));
 NOR3_X4 _04388_ (.A1(_00697_),
    .A2(net12),
    .A3(net13),
    .ZN(_00708_));
 NAND2_X4 _04389_ (.A1(_00675_),
    .A2(_00708_),
    .ZN(_00709_));
 NOR2_X1 _04390_ (.A1(_00656_),
    .A2(_00709_),
    .ZN(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__20.cg_i.en_i ));
 NOR3_X4 _04391_ (.A1(_00697_),
    .A2(_00666_),
    .A3(net13),
    .ZN(_00710_));
 NAND2_X4 _04392_ (.A1(_00675_),
    .A2(_00710_),
    .ZN(_00711_));
 NOR2_X1 _04393_ (.A1(_00656_),
    .A2(_00711_),
    .ZN(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__21.cg_i.en_i ));
 NAND2_X4 _04394_ (.A1(_00675_),
    .A2(_00701_),
    .ZN(_00712_));
 NOR2_X1 _04395_ (.A1(_00656_),
    .A2(_00712_),
    .ZN(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__22.cg_i.en_i ));
 NAND2_X4 _04396_ (.A1(_00675_),
    .A2(_00705_),
    .ZN(_00713_));
 NOR2_X1 _04397_ (.A1(_00656_),
    .A2(_00713_),
    .ZN(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__23.cg_i.en_i ));
 NAND2_X4 _04398_ (.A1(_00684_),
    .A2(_00708_),
    .ZN(_00714_));
 NOR2_X1 _04399_ (.A1(_00656_),
    .A2(_00714_),
    .ZN(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__24.cg_i.en_i ));
 NAND2_X4 _04400_ (.A1(_00684_),
    .A2(_00710_),
    .ZN(_00715_));
 NOR2_X1 _04401_ (.A1(_00656_),
    .A2(_00715_),
    .ZN(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__25.cg_i.en_i ));
 NAND2_X4 _04402_ (.A1(_00684_),
    .A2(_00701_),
    .ZN(_00716_));
 NOR2_X1 _04403_ (.A1(_00656_),
    .A2(_00716_),
    .ZN(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__26.cg_i.en_i ));
 NAND2_X4 _04404_ (.A1(_00684_),
    .A2(_00705_),
    .ZN(_00717_));
 NOR2_X1 _04405_ (.A1(_00656_),
    .A2(_00717_),
    .ZN(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__27.cg_i.en_i ));
 NAND2_X4 _04406_ (.A1(_00691_),
    .A2(_00708_),
    .ZN(_00718_));
 NOR2_X1 _04407_ (.A1(_00656_),
    .A2(_00718_),
    .ZN(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__28.cg_i.en_i ));
 NAND2_X4 _04408_ (.A1(_00691_),
    .A2(_00710_),
    .ZN(_00719_));
 NOR2_X1 _04409_ (.A1(_00656_),
    .A2(_00719_),
    .ZN(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__29.cg_i.en_i ));
 NAND2_X4 _04410_ (.A1(_00691_),
    .A2(_00701_),
    .ZN(_00720_));
 NOR2_X1 _04411_ (.A1(_00656_),
    .A2(_00720_),
    .ZN(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__30.cg_i.en_i ));
 NAND2_X4 _04412_ (.A1(_00691_),
    .A2(_00705_),
    .ZN(_00721_));
 NOR2_X1 _04413_ (.A1(_00656_),
    .A2(_00721_),
    .ZN(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__31.cg_i.en_i ));
 INV_X1 _04414_ (.A(net18),
    .ZN(_00722_));
 NOR2_X4 _04415_ (.A1(_00722_),
    .A2(net17),
    .ZN(_00723_));
 NAND2_X4 _04416_ (.A1(_00655_),
    .A2(_00723_),
    .ZN(_00724_));
 BUF_X8 max_cap214 (.A(net216),
    .Z(net214));
 INV_X1 _04418_ (.A(_00724_),
    .ZN(\lut.gen_sub_units_scm.__14.sub_unit_i.cg_we_global.en_i ));
 BUF_X8 max_cap213 (.A(net214),
    .Z(net213));
 NOR2_X1 _04420_ (.A1(_00665_),
    .A2(_00724_),
    .ZN(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__0.cg_i.en_i ));
 BUF_X4 max_cap212 (.A(_01002_),
    .Z(net212));
 NOR2_X1 _04422_ (.A1(_00668_),
    .A2(_00724_),
    .ZN(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__1.cg_i.en_i ));
 BUF_X8 max_cap211 (.A(net212),
    .Z(net211));
 NOR2_X1 _04424_ (.A1(_00671_),
    .A2(_00724_),
    .ZN(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__2.cg_i.en_i ));
 BUF_X4 max_cap210 (.A(net212),
    .Z(net210));
 NOR2_X1 _04426_ (.A1(_00673_),
    .A2(_00724_),
    .ZN(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__3.cg_i.en_i ));
 BUF_X8 max_cap209 (.A(net210),
    .Z(net209));
 NOR2_X1 _04428_ (.A1(_00678_),
    .A2(_00724_),
    .ZN(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__4.cg_i.en_i ));
 BUF_X4 wire208 (.A(net212),
    .Z(net208));
 NOR2_X1 _04430_ (.A1(_00680_),
    .A2(_00724_),
    .ZN(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__5.cg_i.en_i ));
 BUF_X4 max_cap207 (.A(net211),
    .Z(net207));
 NOR2_X1 _04432_ (.A1(_00681_),
    .A2(_00724_),
    .ZN(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__6.cg_i.en_i ));
 BUF_X16 max_cap206 (.A(_01007_),
    .Z(net206));
 NOR2_X1 _04434_ (.A1(_00682_),
    .A2(_00724_),
    .ZN(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__7.cg_i.en_i ));
 BUF_X16 max_cap205 (.A(_01007_),
    .Z(net205));
 NOR2_X1 _04436_ (.A1(_00686_),
    .A2(_00724_),
    .ZN(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__8.cg_i.en_i ));
 BUF_X16 max_cap204 (.A(net205),
    .Z(net204));
 BUF_X16 max_cap203 (.A(_01007_),
    .Z(net203));
 NOR2_X1 _04439_ (.A1(_00688_),
    .A2(_00724_),
    .ZN(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__9.cg_i.en_i ));
 BUF_X8 max_cap202 (.A(_01009_),
    .Z(net202));
 NOR2_X1 _04441_ (.A1(_00689_),
    .A2(_00724_),
    .ZN(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__10.cg_i.en_i ));
 BUF_X8 max_cap201 (.A(net202),
    .Z(net201));
 NOR2_X1 _04443_ (.A1(_00690_),
    .A2(_00724_),
    .ZN(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__11.cg_i.en_i ));
 BUF_X8 max_cap200 (.A(net201),
    .Z(net200));
 NOR2_X1 _04445_ (.A1(_00693_),
    .A2(_00724_),
    .ZN(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__12.cg_i.en_i ));
 BUF_X4 max_cap199 (.A(net202),
    .Z(net199));
 NOR2_X1 _04447_ (.A1(_00694_),
    .A2(_00724_),
    .ZN(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__13.cg_i.en_i ));
 BUF_X8 max_cap198 (.A(_01009_),
    .Z(net198));
 NOR2_X1 _04449_ (.A1(_00695_),
    .A2(_00724_),
    .ZN(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__14.cg_i.en_i ));
 BUF_X4 wire197 (.A(net198),
    .Z(net197));
 NOR2_X1 _04451_ (.A1(_00696_),
    .A2(_00724_),
    .ZN(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__15.cg_i.en_i ));
 BUF_X4 wire196 (.A(_01009_),
    .Z(net196));
 NOR2_X1 _04453_ (.A1(_00699_),
    .A2(_00724_),
    .ZN(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__16.cg_i.en_i ));
 BUF_X8 max_cap195 (.A(net196),
    .Z(net195));
 NOR2_X1 _04455_ (.A1(_00700_),
    .A2(_00724_),
    .ZN(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__17.cg_i.en_i ));
 BUF_X8 max_cap194 (.A(net195),
    .Z(net194));
 NOR2_X1 _04457_ (.A1(_00703_),
    .A2(_00724_),
    .ZN(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__18.cg_i.en_i ));
 BUF_X4 max_cap193 (.A(net196),
    .Z(net193));
 BUF_X8 max_cap192 (.A(_01021_),
    .Z(net192));
 NOR2_X1 _04460_ (.A1(_00707_),
    .A2(_00724_),
    .ZN(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__19.cg_i.en_i ));
 BUF_X8 max_cap191 (.A(net192),
    .Z(net191));
 NOR2_X1 _04462_ (.A1(_00709_),
    .A2(_00724_),
    .ZN(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__20.cg_i.en_i ));
 BUF_X8 wire190 (.A(net191),
    .Z(net190));
 NOR2_X1 _04464_ (.A1(_00711_),
    .A2(_00724_),
    .ZN(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__21.cg_i.en_i ));
 BUF_X16 max_cap189 (.A(net190),
    .Z(net189));
 NOR2_X1 _04466_ (.A1(_00712_),
    .A2(_00724_),
    .ZN(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__22.cg_i.en_i ));
 BUF_X8 max_cap188 (.A(net192),
    .Z(net188));
 NOR2_X1 _04468_ (.A1(_00713_),
    .A2(_00724_),
    .ZN(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__23.cg_i.en_i ));
 BUF_X8 max_cap187 (.A(_01021_),
    .Z(net187));
 NOR2_X1 _04470_ (.A1(_00714_),
    .A2(_00724_),
    .ZN(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__24.cg_i.en_i ));
 BUF_X8 max_cap186 (.A(net187),
    .Z(net186));
 NOR2_X1 _04472_ (.A1(_00715_),
    .A2(_00724_),
    .ZN(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__25.cg_i.en_i ));
 BUF_X8 max_cap185 (.A(_01034_),
    .Z(net185));
 NOR2_X1 _04474_ (.A1(_00716_),
    .A2(_00724_),
    .ZN(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__26.cg_i.en_i ));
 BUF_X4 wire184 (.A(_01034_),
    .Z(net184));
 NOR2_X1 _04476_ (.A1(_00717_),
    .A2(_00724_),
    .ZN(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__27.cg_i.en_i ));
 BUF_X4 max_cap183 (.A(_01034_),
    .Z(net183));
 NOR2_X1 _04478_ (.A1(_00718_),
    .A2(_00724_),
    .ZN(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__28.cg_i.en_i ));
 BUF_X4 max_cap182 (.A(net183),
    .Z(net182));
 NOR2_X1 _04480_ (.A1(_00719_),
    .A2(_00724_),
    .ZN(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__29.cg_i.en_i ));
 BUF_X4 max_cap181 (.A(_01034_),
    .Z(net181));
 NOR2_X1 _04482_ (.A1(_00720_),
    .A2(_00724_),
    .ZN(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__30.cg_i.en_i ));
 BUF_X8 max_cap180 (.A(net181),
    .Z(net180));
 NOR2_X1 _04484_ (.A1(_00721_),
    .A2(_00724_),
    .ZN(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__31.cg_i.en_i ));
 AND2_X4 _04485_ (.A1(_00722_),
    .A2(net17),
    .ZN(_00760_));
 NAND2_X4 _04486_ (.A1(_00655_),
    .A2(_00760_),
    .ZN(_00761_));
 BUF_X4 max_cap179 (.A(net181),
    .Z(net179));
 INV_X1 _04488_ (.A(_00761_),
    .ZN(\lut.gen_sub_units_scm.__13.sub_unit_i.cg_we_global.en_i ));
 NOR2_X1 _04489_ (.A1(_00665_),
    .A2(_00761_),
    .ZN(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__0.cg_i.en_i ));
 NOR2_X1 _04490_ (.A1(_00668_),
    .A2(_00761_),
    .ZN(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__1.cg_i.en_i ));
 NOR2_X1 _04491_ (.A1(_00671_),
    .A2(_00761_),
    .ZN(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__2.cg_i.en_i ));
 NOR2_X1 _04492_ (.A1(_00673_),
    .A2(_00761_),
    .ZN(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__3.cg_i.en_i ));
 NOR2_X1 _04493_ (.A1(_00678_),
    .A2(_00761_),
    .ZN(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__4.cg_i.en_i ));
 NOR2_X1 _04494_ (.A1(_00680_),
    .A2(_00761_),
    .ZN(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__5.cg_i.en_i ));
 NOR2_X1 _04495_ (.A1(_00681_),
    .A2(_00761_),
    .ZN(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__6.cg_i.en_i ));
 NOR2_X1 _04496_ (.A1(_00682_),
    .A2(_00761_),
    .ZN(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__7.cg_i.en_i ));
 NOR2_X1 _04497_ (.A1(_00686_),
    .A2(_00761_),
    .ZN(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__8.cg_i.en_i ));
 BUF_X4 max_cap178 (.A(net180),
    .Z(net178));
 NOR2_X1 _04499_ (.A1(_00688_),
    .A2(_00761_),
    .ZN(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__9.cg_i.en_i ));
 NOR2_X1 _04500_ (.A1(_00689_),
    .A2(_00761_),
    .ZN(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__10.cg_i.en_i ));
 NOR2_X1 _04501_ (.A1(_00690_),
    .A2(_00761_),
    .ZN(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__11.cg_i.en_i ));
 NOR2_X1 _04502_ (.A1(_00693_),
    .A2(_00761_),
    .ZN(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__12.cg_i.en_i ));
 NOR2_X1 _04503_ (.A1(_00694_),
    .A2(_00761_),
    .ZN(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__13.cg_i.en_i ));
 NOR2_X1 _04504_ (.A1(_00695_),
    .A2(_00761_),
    .ZN(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__14.cg_i.en_i ));
 NOR2_X1 _04505_ (.A1(_00696_),
    .A2(_00761_),
    .ZN(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__15.cg_i.en_i ));
 NOR2_X1 _04506_ (.A1(_00699_),
    .A2(_00761_),
    .ZN(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__16.cg_i.en_i ));
 NOR2_X1 _04507_ (.A1(_00700_),
    .A2(_00761_),
    .ZN(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__17.cg_i.en_i ));
 NOR2_X1 _04508_ (.A1(_00703_),
    .A2(_00761_),
    .ZN(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__18.cg_i.en_i ));
 BUF_X8 max_cap177 (.A(net185),
    .Z(net177));
 NOR2_X1 _04510_ (.A1(_00707_),
    .A2(_00761_),
    .ZN(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__19.cg_i.en_i ));
 NOR2_X1 _04511_ (.A1(_00709_),
    .A2(_00761_),
    .ZN(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__20.cg_i.en_i ));
 NOR2_X1 _04512_ (.A1(_00711_),
    .A2(_00761_),
    .ZN(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__21.cg_i.en_i ));
 NOR2_X1 _04513_ (.A1(_00712_),
    .A2(_00761_),
    .ZN(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__22.cg_i.en_i ));
 NOR2_X1 _04514_ (.A1(_00713_),
    .A2(_00761_),
    .ZN(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__23.cg_i.en_i ));
 NOR2_X1 _04515_ (.A1(_00714_),
    .A2(_00761_),
    .ZN(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__24.cg_i.en_i ));
 NOR2_X1 _04516_ (.A1(_00715_),
    .A2(_00761_),
    .ZN(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__25.cg_i.en_i ));
 NOR2_X1 _04517_ (.A1(_00716_),
    .A2(_00761_),
    .ZN(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__26.cg_i.en_i ));
 NOR2_X1 _04518_ (.A1(_00717_),
    .A2(_00761_),
    .ZN(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__27.cg_i.en_i ));
 NOR2_X1 _04519_ (.A1(_00718_),
    .A2(_00761_),
    .ZN(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__28.cg_i.en_i ));
 NOR2_X1 _04520_ (.A1(_00719_),
    .A2(_00761_),
    .ZN(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__29.cg_i.en_i ));
 NOR2_X1 _04521_ (.A1(_00720_),
    .A2(_00761_),
    .ZN(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__30.cg_i.en_i ));
 NOR2_X1 _04522_ (.A1(_00721_),
    .A2(_00761_),
    .ZN(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__31.cg_i.en_i ));
 NOR2_X4 _04523_ (.A1(net18),
    .A2(net17),
    .ZN(_00765_));
 NAND2_X4 _04524_ (.A1(_00655_),
    .A2(_00765_),
    .ZN(_00766_));
 BUF_X8 max_cap176 (.A(net177),
    .Z(net176));
 INV_X1 _04526_ (.A(_00766_),
    .ZN(\lut.gen_sub_units_scm.__12.sub_unit_i.cg_we_global.en_i ));
 NOR2_X1 _04527_ (.A1(_00665_),
    .A2(_00766_),
    .ZN(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__0.cg_i.en_i ));
 NOR2_X1 _04528_ (.A1(_00668_),
    .A2(_00766_),
    .ZN(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__1.cg_i.en_i ));
 NOR2_X1 _04529_ (.A1(_00671_),
    .A2(_00766_),
    .ZN(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__2.cg_i.en_i ));
 NOR2_X1 _04530_ (.A1(_00673_),
    .A2(_00766_),
    .ZN(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__3.cg_i.en_i ));
 NOR2_X1 _04531_ (.A1(_00678_),
    .A2(_00766_),
    .ZN(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__4.cg_i.en_i ));
 NOR2_X1 _04532_ (.A1(_00680_),
    .A2(_00766_),
    .ZN(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__5.cg_i.en_i ));
 NOR2_X1 _04533_ (.A1(_00681_),
    .A2(_00766_),
    .ZN(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__6.cg_i.en_i ));
 NOR2_X1 _04534_ (.A1(_00682_),
    .A2(_00766_),
    .ZN(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__7.cg_i.en_i ));
 NOR2_X1 _04535_ (.A1(_00686_),
    .A2(_00766_),
    .ZN(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__8.cg_i.en_i ));
 BUF_X4 max_cap175 (.A(_01038_),
    .Z(net175));
 NOR2_X1 _04537_ (.A1(_00688_),
    .A2(_00766_),
    .ZN(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__9.cg_i.en_i ));
 NOR2_X1 _04538_ (.A1(_00689_),
    .A2(_00766_),
    .ZN(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__10.cg_i.en_i ));
 NOR2_X1 _04539_ (.A1(_00690_),
    .A2(_00766_),
    .ZN(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__11.cg_i.en_i ));
 NOR2_X1 _04540_ (.A1(_00693_),
    .A2(_00766_),
    .ZN(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__12.cg_i.en_i ));
 NOR2_X1 _04541_ (.A1(_00694_),
    .A2(_00766_),
    .ZN(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__13.cg_i.en_i ));
 NOR2_X1 _04542_ (.A1(_00695_),
    .A2(_00766_),
    .ZN(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__14.cg_i.en_i ));
 NOR2_X1 _04543_ (.A1(_00696_),
    .A2(_00766_),
    .ZN(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__15.cg_i.en_i ));
 NOR2_X1 _04544_ (.A1(_00699_),
    .A2(_00766_),
    .ZN(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__16.cg_i.en_i ));
 NOR2_X1 _04545_ (.A1(_00700_),
    .A2(_00766_),
    .ZN(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__17.cg_i.en_i ));
 NOR2_X1 _04546_ (.A1(_00703_),
    .A2(_00766_),
    .ZN(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__18.cg_i.en_i ));
 BUF_X8 max_cap174 (.A(net175),
    .Z(net174));
 NOR2_X1 _04548_ (.A1(_00707_),
    .A2(_00766_),
    .ZN(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__19.cg_i.en_i ));
 NOR2_X1 _04549_ (.A1(_00709_),
    .A2(_00766_),
    .ZN(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__20.cg_i.en_i ));
 NOR2_X1 _04550_ (.A1(_00711_),
    .A2(_00766_),
    .ZN(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__21.cg_i.en_i ));
 NOR2_X1 _04551_ (.A1(_00712_),
    .A2(_00766_),
    .ZN(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__22.cg_i.en_i ));
 NOR2_X1 _04552_ (.A1(_00713_),
    .A2(_00766_),
    .ZN(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__23.cg_i.en_i ));
 NOR2_X1 _04553_ (.A1(_00714_),
    .A2(_00766_),
    .ZN(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__24.cg_i.en_i ));
 NOR2_X1 _04554_ (.A1(_00715_),
    .A2(_00766_),
    .ZN(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__25.cg_i.en_i ));
 NOR2_X1 _04555_ (.A1(_00716_),
    .A2(_00766_),
    .ZN(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__26.cg_i.en_i ));
 NOR2_X1 _04556_ (.A1(_00717_),
    .A2(_00766_),
    .ZN(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__27.cg_i.en_i ));
 NOR2_X1 _04557_ (.A1(_00718_),
    .A2(_00766_),
    .ZN(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__28.cg_i.en_i ));
 NOR2_X1 _04558_ (.A1(_00719_),
    .A2(_00766_),
    .ZN(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__29.cg_i.en_i ));
 NOR2_X1 _04559_ (.A1(_00720_),
    .A2(_00766_),
    .ZN(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__30.cg_i.en_i ));
 NOR2_X1 _04560_ (.A1(_00721_),
    .A2(_00766_),
    .ZN(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__31.cg_i.en_i ));
 INV_X1 _04561_ (.A(net19),
    .ZN(_00770_));
 AND3_X4 _04562_ (.A1(net20),
    .A2(_00770_),
    .A3(net29),
    .ZN(_00771_));
 BUF_X8 max_cap173 (.A(net175),
    .Z(net173));
 NAND3_X4 _04564_ (.A1(net18),
    .A2(net17),
    .A3(_00771_),
    .ZN(_00773_));
 BUF_X4 max_cap172 (.A(_01038_),
    .Z(net172));
 INV_X1 _04566_ (.A(_00773_),
    .ZN(\lut.gen_sub_units_scm.__11.sub_unit_i.cg_we_global.en_i ));
 NOR2_X1 _04567_ (.A1(_00665_),
    .A2(_00773_),
    .ZN(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__0.cg_i.en_i ));
 NOR2_X1 _04568_ (.A1(_00668_),
    .A2(_00773_),
    .ZN(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__1.cg_i.en_i ));
 NOR2_X1 _04569_ (.A1(_00671_),
    .A2(_00773_),
    .ZN(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__2.cg_i.en_i ));
 NOR2_X1 _04570_ (.A1(_00673_),
    .A2(_00773_),
    .ZN(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__3.cg_i.en_i ));
 NOR2_X1 _04571_ (.A1(_00678_),
    .A2(_00773_),
    .ZN(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__4.cg_i.en_i ));
 NOR2_X1 _04572_ (.A1(_00680_),
    .A2(_00773_),
    .ZN(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__5.cg_i.en_i ));
 NOR2_X1 _04573_ (.A1(_00681_),
    .A2(_00773_),
    .ZN(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__6.cg_i.en_i ));
 NOR2_X1 _04574_ (.A1(_00682_),
    .A2(_00773_),
    .ZN(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__7.cg_i.en_i ));
 NOR2_X1 _04575_ (.A1(_00686_),
    .A2(_00773_),
    .ZN(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__8.cg_i.en_i ));
 BUF_X4 max_cap171 (.A(_01038_),
    .Z(net171));
 NOR2_X1 _04577_ (.A1(_00688_),
    .A2(_00773_),
    .ZN(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__9.cg_i.en_i ));
 NOR2_X1 _04578_ (.A1(_00689_),
    .A2(_00773_),
    .ZN(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__10.cg_i.en_i ));
 NOR2_X1 _04579_ (.A1(_00690_),
    .A2(_00773_),
    .ZN(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__11.cg_i.en_i ));
 NOR2_X1 _04580_ (.A1(_00693_),
    .A2(_00773_),
    .ZN(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__12.cg_i.en_i ));
 NOR2_X1 _04581_ (.A1(_00694_),
    .A2(_00773_),
    .ZN(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__13.cg_i.en_i ));
 NOR2_X1 _04582_ (.A1(_00695_),
    .A2(_00773_),
    .ZN(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__14.cg_i.en_i ));
 NOR2_X1 _04583_ (.A1(_00696_),
    .A2(_00773_),
    .ZN(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__15.cg_i.en_i ));
 NOR2_X1 _04584_ (.A1(_00699_),
    .A2(_00773_),
    .ZN(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__16.cg_i.en_i ));
 NOR2_X1 _04585_ (.A1(_00700_),
    .A2(_00773_),
    .ZN(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__17.cg_i.en_i ));
 NOR2_X1 _04586_ (.A1(_00703_),
    .A2(_00773_),
    .ZN(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__18.cg_i.en_i ));
 BUF_X4 max_cap170 (.A(_01038_),
    .Z(net170));
 NOR2_X1 _04588_ (.A1(_00707_),
    .A2(_00773_),
    .ZN(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__19.cg_i.en_i ));
 NOR2_X1 _04589_ (.A1(_00709_),
    .A2(_00773_),
    .ZN(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__20.cg_i.en_i ));
 NOR2_X1 _04590_ (.A1(_00711_),
    .A2(_00773_),
    .ZN(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__21.cg_i.en_i ));
 NOR2_X1 _04591_ (.A1(_00712_),
    .A2(_00773_),
    .ZN(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__22.cg_i.en_i ));
 NOR2_X1 _04592_ (.A1(_00713_),
    .A2(_00773_),
    .ZN(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__23.cg_i.en_i ));
 NOR2_X1 _04593_ (.A1(_00714_),
    .A2(_00773_),
    .ZN(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__24.cg_i.en_i ));
 NOR2_X1 _04594_ (.A1(_00715_),
    .A2(_00773_),
    .ZN(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__25.cg_i.en_i ));
 NOR2_X1 _04595_ (.A1(_00716_),
    .A2(_00773_),
    .ZN(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__26.cg_i.en_i ));
 NOR2_X1 _04596_ (.A1(_00717_),
    .A2(_00773_),
    .ZN(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__27.cg_i.en_i ));
 NOR2_X1 _04597_ (.A1(_00718_),
    .A2(_00773_),
    .ZN(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__28.cg_i.en_i ));
 NOR2_X1 _04598_ (.A1(_00719_),
    .A2(_00773_),
    .ZN(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__29.cg_i.en_i ));
 NOR2_X1 _04599_ (.A1(_00720_),
    .A2(_00773_),
    .ZN(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__30.cg_i.en_i ));
 NOR2_X1 _04600_ (.A1(_00721_),
    .A2(_00773_),
    .ZN(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__31.cg_i.en_i ));
 NAND2_X4 _04601_ (.A1(_00723_),
    .A2(_00771_),
    .ZN(_00777_));
 BUF_X8 max_cap169 (.A(net170),
    .Z(net169));
 INV_X1 _04603_ (.A(_00777_),
    .ZN(\lut.gen_sub_units_scm.__10.sub_unit_i.cg_we_global.en_i ));
 NOR2_X1 _04604_ (.A1(_00665_),
    .A2(_00777_),
    .ZN(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__0.cg_i.en_i ));
 NOR2_X1 _04605_ (.A1(_00668_),
    .A2(_00777_),
    .ZN(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__1.cg_i.en_i ));
 NOR2_X1 _04606_ (.A1(_00671_),
    .A2(_00777_),
    .ZN(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__2.cg_i.en_i ));
 NOR2_X1 _04607_ (.A1(_00673_),
    .A2(_00777_),
    .ZN(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__3.cg_i.en_i ));
 NOR2_X1 _04608_ (.A1(_00678_),
    .A2(_00777_),
    .ZN(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__4.cg_i.en_i ));
 NOR2_X1 _04609_ (.A1(_00680_),
    .A2(_00777_),
    .ZN(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__5.cg_i.en_i ));
 NOR2_X1 _04610_ (.A1(_00681_),
    .A2(_00777_),
    .ZN(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__6.cg_i.en_i ));
 NOR2_X1 _04611_ (.A1(_00682_),
    .A2(_00777_),
    .ZN(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__7.cg_i.en_i ));
 NOR2_X1 _04612_ (.A1(_00686_),
    .A2(_00777_),
    .ZN(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__8.cg_i.en_i ));
 BUF_X4 wire168 (.A(_01038_),
    .Z(net168));
 NOR2_X1 _04614_ (.A1(_00688_),
    .A2(_00777_),
    .ZN(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__9.cg_i.en_i ));
 NOR2_X1 _04615_ (.A1(_00689_),
    .A2(_00777_),
    .ZN(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__10.cg_i.en_i ));
 NOR2_X1 _04616_ (.A1(_00690_),
    .A2(_00777_),
    .ZN(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__11.cg_i.en_i ));
 NOR2_X1 _04617_ (.A1(_00693_),
    .A2(_00777_),
    .ZN(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__12.cg_i.en_i ));
 NOR2_X1 _04618_ (.A1(_00694_),
    .A2(_00777_),
    .ZN(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__13.cg_i.en_i ));
 NOR2_X1 _04619_ (.A1(_00695_),
    .A2(_00777_),
    .ZN(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__14.cg_i.en_i ));
 NOR2_X1 _04620_ (.A1(_00696_),
    .A2(_00777_),
    .ZN(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__15.cg_i.en_i ));
 NOR2_X1 _04621_ (.A1(_00699_),
    .A2(_00777_),
    .ZN(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__16.cg_i.en_i ));
 NOR2_X1 _04622_ (.A1(_00700_),
    .A2(_00777_),
    .ZN(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__17.cg_i.en_i ));
 NOR2_X1 _04623_ (.A1(_00703_),
    .A2(_00777_),
    .ZN(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__18.cg_i.en_i ));
 BUF_X4 max_cap167 (.A(net172),
    .Z(net167));
 NOR2_X1 _04625_ (.A1(_00707_),
    .A2(_00777_),
    .ZN(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__19.cg_i.en_i ));
 NOR2_X1 _04626_ (.A1(_00709_),
    .A2(_00777_),
    .ZN(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__20.cg_i.en_i ));
 NOR2_X1 _04627_ (.A1(_00711_),
    .A2(_00777_),
    .ZN(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__21.cg_i.en_i ));
 NOR2_X1 _04628_ (.A1(_00712_),
    .A2(_00777_),
    .ZN(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__22.cg_i.en_i ));
 NOR2_X1 _04629_ (.A1(_00713_),
    .A2(_00777_),
    .ZN(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__23.cg_i.en_i ));
 NOR2_X1 _04630_ (.A1(_00714_),
    .A2(_00777_),
    .ZN(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__24.cg_i.en_i ));
 NOR2_X1 _04631_ (.A1(_00715_),
    .A2(_00777_),
    .ZN(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__25.cg_i.en_i ));
 NOR2_X1 _04632_ (.A1(_00716_),
    .A2(_00777_),
    .ZN(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__26.cg_i.en_i ));
 NOR2_X1 _04633_ (.A1(_00717_),
    .A2(_00777_),
    .ZN(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__27.cg_i.en_i ));
 NOR2_X1 _04634_ (.A1(_00718_),
    .A2(_00777_),
    .ZN(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__28.cg_i.en_i ));
 NOR2_X1 _04635_ (.A1(_00719_),
    .A2(_00777_),
    .ZN(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__29.cg_i.en_i ));
 NOR2_X1 _04636_ (.A1(_00720_),
    .A2(_00777_),
    .ZN(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__30.cg_i.en_i ));
 NOR2_X1 _04637_ (.A1(_00721_),
    .A2(_00777_),
    .ZN(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__31.cg_i.en_i ));
 NAND2_X4 _04638_ (.A1(_00760_),
    .A2(_00771_),
    .ZN(_00781_));
 BUF_X8 max_cap166 (.A(net167),
    .Z(net166));
 INV_X1 _04640_ (.A(_00781_),
    .ZN(\lut.gen_sub_units_scm.__9.sub_unit_i.cg_we_global.en_i ));
 NOR2_X1 _04641_ (.A1(_00665_),
    .A2(_00781_),
    .ZN(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__0.cg_i.en_i ));
 NOR2_X1 _04642_ (.A1(_00668_),
    .A2(_00781_),
    .ZN(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__1.cg_i.en_i ));
 NOR2_X1 _04643_ (.A1(_00671_),
    .A2(_00781_),
    .ZN(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__2.cg_i.en_i ));
 NOR2_X1 _04644_ (.A1(_00673_),
    .A2(_00781_),
    .ZN(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__3.cg_i.en_i ));
 NOR2_X1 _04645_ (.A1(_00678_),
    .A2(_00781_),
    .ZN(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__4.cg_i.en_i ));
 NOR2_X1 _04646_ (.A1(_00680_),
    .A2(_00781_),
    .ZN(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__5.cg_i.en_i ));
 NOR2_X1 _04647_ (.A1(_00681_),
    .A2(_00781_),
    .ZN(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__6.cg_i.en_i ));
 NOR2_X1 _04648_ (.A1(_00682_),
    .A2(_00781_),
    .ZN(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__7.cg_i.en_i ));
 NOR2_X1 _04649_ (.A1(_00686_),
    .A2(_00781_),
    .ZN(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__8.cg_i.en_i ));
 BUF_X4 max_cap165 (.A(_01042_),
    .Z(net165));
 NOR2_X1 _04651_ (.A1(_00688_),
    .A2(_00781_),
    .ZN(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__9.cg_i.en_i ));
 NOR2_X1 _04652_ (.A1(_00689_),
    .A2(_00781_),
    .ZN(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__10.cg_i.en_i ));
 NOR2_X1 _04653_ (.A1(_00690_),
    .A2(_00781_),
    .ZN(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__11.cg_i.en_i ));
 NOR2_X1 _04654_ (.A1(_00693_),
    .A2(_00781_),
    .ZN(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__12.cg_i.en_i ));
 NOR2_X1 _04655_ (.A1(_00694_),
    .A2(_00781_),
    .ZN(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__13.cg_i.en_i ));
 NOR2_X1 _04656_ (.A1(_00695_),
    .A2(_00781_),
    .ZN(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__14.cg_i.en_i ));
 NOR2_X1 _04657_ (.A1(_00696_),
    .A2(_00781_),
    .ZN(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__15.cg_i.en_i ));
 NOR2_X1 _04658_ (.A1(_00699_),
    .A2(_00781_),
    .ZN(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__16.cg_i.en_i ));
 NOR2_X1 _04659_ (.A1(_00700_),
    .A2(_00781_),
    .ZN(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__17.cg_i.en_i ));
 NOR2_X1 _04660_ (.A1(_00703_),
    .A2(_00781_),
    .ZN(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__18.cg_i.en_i ));
 BUF_X8 max_cap164 (.A(_01042_),
    .Z(net164));
 NOR2_X1 _04662_ (.A1(_00707_),
    .A2(_00781_),
    .ZN(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__19.cg_i.en_i ));
 NOR2_X1 _04663_ (.A1(_00709_),
    .A2(_00781_),
    .ZN(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__20.cg_i.en_i ));
 NOR2_X1 _04664_ (.A1(_00711_),
    .A2(_00781_),
    .ZN(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__21.cg_i.en_i ));
 NOR2_X1 _04665_ (.A1(_00712_),
    .A2(_00781_),
    .ZN(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__22.cg_i.en_i ));
 NOR2_X1 _04666_ (.A1(_00713_),
    .A2(_00781_),
    .ZN(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__23.cg_i.en_i ));
 NOR2_X1 _04667_ (.A1(_00714_),
    .A2(_00781_),
    .ZN(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__24.cg_i.en_i ));
 NOR2_X1 _04668_ (.A1(_00715_),
    .A2(_00781_),
    .ZN(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__25.cg_i.en_i ));
 NOR2_X1 _04669_ (.A1(_00716_),
    .A2(_00781_),
    .ZN(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__26.cg_i.en_i ));
 NOR2_X1 _04670_ (.A1(_00717_),
    .A2(_00781_),
    .ZN(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__27.cg_i.en_i ));
 NOR2_X1 _04671_ (.A1(_00718_),
    .A2(_00781_),
    .ZN(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__28.cg_i.en_i ));
 NOR2_X1 _04672_ (.A1(_00719_),
    .A2(_00781_),
    .ZN(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__29.cg_i.en_i ));
 NOR2_X1 _04673_ (.A1(_00720_),
    .A2(_00781_),
    .ZN(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__30.cg_i.en_i ));
 NOR2_X1 _04674_ (.A1(_00721_),
    .A2(_00781_),
    .ZN(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__31.cg_i.en_i ));
 NAND2_X4 _04675_ (.A1(_00765_),
    .A2(_00771_),
    .ZN(_00785_));
 BUF_X4 wire163 (.A(net164),
    .Z(net163));
 INV_X1 _04677_ (.A(_00785_),
    .ZN(\lut.gen_sub_units_scm.__8.sub_unit_i.cg_we_global.en_i ));
 NOR2_X1 _04678_ (.A1(_00665_),
    .A2(_00785_),
    .ZN(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__0.cg_i.en_i ));
 NOR2_X1 _04679_ (.A1(_00668_),
    .A2(_00785_),
    .ZN(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__1.cg_i.en_i ));
 NOR2_X1 _04680_ (.A1(_00671_),
    .A2(_00785_),
    .ZN(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__2.cg_i.en_i ));
 NOR2_X1 _04681_ (.A1(_00673_),
    .A2(_00785_),
    .ZN(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__3.cg_i.en_i ));
 NOR2_X1 _04682_ (.A1(_00678_),
    .A2(_00785_),
    .ZN(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__4.cg_i.en_i ));
 NOR2_X1 _04683_ (.A1(_00680_),
    .A2(_00785_),
    .ZN(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__5.cg_i.en_i ));
 NOR2_X1 _04684_ (.A1(_00681_),
    .A2(_00785_),
    .ZN(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__6.cg_i.en_i ));
 NOR2_X1 _04685_ (.A1(_00682_),
    .A2(_00785_),
    .ZN(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__7.cg_i.en_i ));
 NOR2_X1 _04686_ (.A1(_00686_),
    .A2(_00785_),
    .ZN(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__8.cg_i.en_i ));
 BUF_X4 max_cap162 (.A(net163),
    .Z(net162));
 NOR2_X1 _04688_ (.A1(_00688_),
    .A2(_00785_),
    .ZN(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__9.cg_i.en_i ));
 NOR2_X1 _04689_ (.A1(_00689_),
    .A2(_00785_),
    .ZN(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__10.cg_i.en_i ));
 NOR2_X1 _04690_ (.A1(_00690_),
    .A2(_00785_),
    .ZN(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__11.cg_i.en_i ));
 NOR2_X1 _04691_ (.A1(_00693_),
    .A2(_00785_),
    .ZN(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__12.cg_i.en_i ));
 NOR2_X1 _04692_ (.A1(_00694_),
    .A2(_00785_),
    .ZN(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__13.cg_i.en_i ));
 NOR2_X1 _04693_ (.A1(_00695_),
    .A2(_00785_),
    .ZN(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__14.cg_i.en_i ));
 NOR2_X1 _04694_ (.A1(_00696_),
    .A2(_00785_),
    .ZN(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__15.cg_i.en_i ));
 NOR2_X1 _04695_ (.A1(_00699_),
    .A2(_00785_),
    .ZN(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__16.cg_i.en_i ));
 NOR2_X1 _04696_ (.A1(_00700_),
    .A2(_00785_),
    .ZN(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__17.cg_i.en_i ));
 NOR2_X1 _04697_ (.A1(_00703_),
    .A2(_00785_),
    .ZN(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__18.cg_i.en_i ));
 BUF_X4 max_cap161 (.A(net164),
    .Z(net161));
 NOR2_X1 _04699_ (.A1(_00707_),
    .A2(_00785_),
    .ZN(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__19.cg_i.en_i ));
 NOR2_X1 _04700_ (.A1(_00709_),
    .A2(_00785_),
    .ZN(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__20.cg_i.en_i ));
 NOR2_X1 _04701_ (.A1(_00711_),
    .A2(_00785_),
    .ZN(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__21.cg_i.en_i ));
 NOR2_X1 _04702_ (.A1(_00712_),
    .A2(_00785_),
    .ZN(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__22.cg_i.en_i ));
 NOR2_X1 _04703_ (.A1(_00713_),
    .A2(_00785_),
    .ZN(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__23.cg_i.en_i ));
 NOR2_X1 _04704_ (.A1(_00714_),
    .A2(_00785_),
    .ZN(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__24.cg_i.en_i ));
 NOR2_X1 _04705_ (.A1(_00715_),
    .A2(_00785_),
    .ZN(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__25.cg_i.en_i ));
 NOR2_X1 _04706_ (.A1(_00716_),
    .A2(_00785_),
    .ZN(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__26.cg_i.en_i ));
 NOR2_X1 _04707_ (.A1(_00717_),
    .A2(_00785_),
    .ZN(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__27.cg_i.en_i ));
 NOR2_X1 _04708_ (.A1(_00718_),
    .A2(_00785_),
    .ZN(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__28.cg_i.en_i ));
 NOR2_X1 _04709_ (.A1(_00719_),
    .A2(_00785_),
    .ZN(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__29.cg_i.en_i ));
 NOR2_X1 _04710_ (.A1(_00720_),
    .A2(_00785_),
    .ZN(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__30.cg_i.en_i ));
 NOR2_X1 _04711_ (.A1(_00721_),
    .A2(_00785_),
    .ZN(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__31.cg_i.en_i ));
 INV_X1 _04712_ (.A(net29),
    .ZN(_00789_));
 NOR3_X4 _04713_ (.A1(net20),
    .A2(_00770_),
    .A3(_00789_),
    .ZN(_00790_));
 NAND3_X4 _04714_ (.A1(net18),
    .A2(net17),
    .A3(_00790_),
    .ZN(_00791_));
 BUF_X4 wire160 (.A(_01042_),
    .Z(net160));
 INV_X1 _04716_ (.A(_00791_),
    .ZN(\lut.gen_sub_units_scm.__7.sub_unit_i.cg_we_global.en_i ));
 NOR2_X1 _04717_ (.A1(_00665_),
    .A2(_00791_),
    .ZN(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__0.cg_i.en_i ));
 NOR2_X1 _04718_ (.A1(_00668_),
    .A2(_00791_),
    .ZN(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__1.cg_i.en_i ));
 NOR2_X1 _04719_ (.A1(_00671_),
    .A2(_00791_),
    .ZN(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__2.cg_i.en_i ));
 NOR2_X1 _04720_ (.A1(_00673_),
    .A2(_00791_),
    .ZN(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__3.cg_i.en_i ));
 NOR2_X1 _04721_ (.A1(_00678_),
    .A2(_00791_),
    .ZN(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__4.cg_i.en_i ));
 NOR2_X1 _04722_ (.A1(_00680_),
    .A2(_00791_),
    .ZN(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__5.cg_i.en_i ));
 NOR2_X1 _04723_ (.A1(_00681_),
    .A2(_00791_),
    .ZN(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__6.cg_i.en_i ));
 NOR2_X1 _04724_ (.A1(_00682_),
    .A2(_00791_),
    .ZN(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__7.cg_i.en_i ));
 NOR2_X1 _04725_ (.A1(_00686_),
    .A2(_00791_),
    .ZN(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__8.cg_i.en_i ));
 BUF_X8 max_cap159 (.A(net165),
    .Z(net159));
 NOR2_X1 _04727_ (.A1(_00688_),
    .A2(_00791_),
    .ZN(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__9.cg_i.en_i ));
 NOR2_X1 _04728_ (.A1(_00689_),
    .A2(_00791_),
    .ZN(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__10.cg_i.en_i ));
 NOR2_X1 _04729_ (.A1(_00690_),
    .A2(_00791_),
    .ZN(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__11.cg_i.en_i ));
 NOR2_X1 _04730_ (.A1(_00693_),
    .A2(_00791_),
    .ZN(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__12.cg_i.en_i ));
 NOR2_X1 _04731_ (.A1(_00694_),
    .A2(_00791_),
    .ZN(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__13.cg_i.en_i ));
 NOR2_X1 _04732_ (.A1(_00695_),
    .A2(_00791_),
    .ZN(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__14.cg_i.en_i ));
 NOR2_X1 _04733_ (.A1(_00696_),
    .A2(_00791_),
    .ZN(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__15.cg_i.en_i ));
 NOR2_X1 _04734_ (.A1(_00699_),
    .A2(_00791_),
    .ZN(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__16.cg_i.en_i ));
 NOR2_X1 _04735_ (.A1(_00700_),
    .A2(_00791_),
    .ZN(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__17.cg_i.en_i ));
 NOR2_X1 _04736_ (.A1(_00703_),
    .A2(_00791_),
    .ZN(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__18.cg_i.en_i ));
 BUF_X4 max_cap158 (.A(net165),
    .Z(net158));
 NOR2_X1 _04738_ (.A1(_00707_),
    .A2(_00791_),
    .ZN(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__19.cg_i.en_i ));
 NOR2_X1 _04739_ (.A1(_00709_),
    .A2(_00791_),
    .ZN(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__20.cg_i.en_i ));
 NOR2_X1 _04740_ (.A1(_00711_),
    .A2(_00791_),
    .ZN(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__21.cg_i.en_i ));
 NOR2_X1 _04741_ (.A1(_00712_),
    .A2(_00791_),
    .ZN(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__22.cg_i.en_i ));
 NOR2_X1 _04742_ (.A1(_00713_),
    .A2(_00791_),
    .ZN(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__23.cg_i.en_i ));
 NOR2_X1 _04743_ (.A1(_00714_),
    .A2(_00791_),
    .ZN(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__24.cg_i.en_i ));
 NOR2_X1 _04744_ (.A1(_00715_),
    .A2(_00791_),
    .ZN(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__25.cg_i.en_i ));
 NOR2_X1 _04745_ (.A1(_00716_),
    .A2(_00791_),
    .ZN(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__26.cg_i.en_i ));
 NOR2_X1 _04746_ (.A1(_00717_),
    .A2(_00791_),
    .ZN(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__27.cg_i.en_i ));
 NOR2_X1 _04747_ (.A1(_00718_),
    .A2(_00791_),
    .ZN(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__28.cg_i.en_i ));
 NOR2_X1 _04748_ (.A1(_00719_),
    .A2(_00791_),
    .ZN(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__29.cg_i.en_i ));
 NOR2_X1 _04749_ (.A1(_00720_),
    .A2(_00791_),
    .ZN(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__30.cg_i.en_i ));
 NOR2_X1 _04750_ (.A1(_00721_),
    .A2(_00791_),
    .ZN(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__31.cg_i.en_i ));
 NAND2_X4 _04751_ (.A1(_00723_),
    .A2(_00790_),
    .ZN(_00795_));
 BUF_X4 max_cap157 (.A(net158),
    .Z(net157));
 INV_X1 _04753_ (.A(_00795_),
    .ZN(\lut.gen_sub_units_scm.__6.sub_unit_i.cg_we_global.en_i ));
 NOR2_X1 _04754_ (.A1(_00665_),
    .A2(_00795_),
    .ZN(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__0.cg_i.en_i ));
 NOR2_X1 _04755_ (.A1(_00668_),
    .A2(_00795_),
    .ZN(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__1.cg_i.en_i ));
 NOR2_X1 _04756_ (.A1(_00671_),
    .A2(_00795_),
    .ZN(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__2.cg_i.en_i ));
 NOR2_X1 _04757_ (.A1(_00673_),
    .A2(_00795_),
    .ZN(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__3.cg_i.en_i ));
 NOR2_X1 _04758_ (.A1(_00678_),
    .A2(_00795_),
    .ZN(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__4.cg_i.en_i ));
 NOR2_X1 _04759_ (.A1(_00680_),
    .A2(_00795_),
    .ZN(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__5.cg_i.en_i ));
 NOR2_X1 _04760_ (.A1(_00681_),
    .A2(_00795_),
    .ZN(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__6.cg_i.en_i ));
 NOR2_X1 _04761_ (.A1(_00682_),
    .A2(_00795_),
    .ZN(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__7.cg_i.en_i ));
 NOR2_X1 _04762_ (.A1(_00686_),
    .A2(_00795_),
    .ZN(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__8.cg_i.en_i ));
 BUF_X8 max_cap156 (.A(net159),
    .Z(net156));
 NOR2_X1 _04764_ (.A1(_00688_),
    .A2(_00795_),
    .ZN(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__9.cg_i.en_i ));
 NOR2_X1 _04765_ (.A1(_00689_),
    .A2(_00795_),
    .ZN(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__10.cg_i.en_i ));
 NOR2_X1 _04766_ (.A1(_00690_),
    .A2(_00795_),
    .ZN(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__11.cg_i.en_i ));
 NOR2_X1 _04767_ (.A1(_00693_),
    .A2(_00795_),
    .ZN(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__12.cg_i.en_i ));
 NOR2_X1 _04768_ (.A1(_00694_),
    .A2(_00795_),
    .ZN(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__13.cg_i.en_i ));
 NOR2_X1 _04769_ (.A1(_00695_),
    .A2(_00795_),
    .ZN(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__14.cg_i.en_i ));
 NOR2_X1 _04770_ (.A1(_00696_),
    .A2(_00795_),
    .ZN(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__15.cg_i.en_i ));
 NOR2_X1 _04771_ (.A1(_00699_),
    .A2(_00795_),
    .ZN(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__16.cg_i.en_i ));
 NOR2_X1 _04772_ (.A1(_00700_),
    .A2(_00795_),
    .ZN(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__17.cg_i.en_i ));
 NOR2_X1 _04773_ (.A1(_00703_),
    .A2(_00795_),
    .ZN(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__18.cg_i.en_i ));
 BUF_X4 max_cap155 (.A(_01046_),
    .Z(net155));
 NOR2_X1 _04775_ (.A1(_00707_),
    .A2(_00795_),
    .ZN(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__19.cg_i.en_i ));
 NOR2_X1 _04776_ (.A1(_00709_),
    .A2(_00795_),
    .ZN(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__20.cg_i.en_i ));
 NOR2_X1 _04777_ (.A1(_00711_),
    .A2(_00795_),
    .ZN(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__21.cg_i.en_i ));
 NOR2_X1 _04778_ (.A1(_00712_),
    .A2(_00795_),
    .ZN(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__22.cg_i.en_i ));
 NOR2_X1 _04779_ (.A1(_00713_),
    .A2(_00795_),
    .ZN(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__23.cg_i.en_i ));
 NOR2_X1 _04780_ (.A1(_00714_),
    .A2(_00795_),
    .ZN(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__24.cg_i.en_i ));
 NOR2_X1 _04781_ (.A1(_00715_),
    .A2(_00795_),
    .ZN(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__25.cg_i.en_i ));
 NOR2_X1 _04782_ (.A1(_00716_),
    .A2(_00795_),
    .ZN(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__26.cg_i.en_i ));
 NOR2_X1 _04783_ (.A1(_00717_),
    .A2(_00795_),
    .ZN(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__27.cg_i.en_i ));
 NOR2_X1 _04784_ (.A1(_00718_),
    .A2(_00795_),
    .ZN(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__28.cg_i.en_i ));
 NOR2_X1 _04785_ (.A1(_00719_),
    .A2(_00795_),
    .ZN(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__29.cg_i.en_i ));
 NOR2_X1 _04786_ (.A1(_00720_),
    .A2(_00795_),
    .ZN(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__30.cg_i.en_i ));
 NOR2_X1 _04787_ (.A1(_00721_),
    .A2(_00795_),
    .ZN(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__31.cg_i.en_i ));
 NAND2_X4 _04788_ (.A1(_00760_),
    .A2(_00790_),
    .ZN(_00799_));
 BUF_X4 max_cap154 (.A(net155),
    .Z(net154));
 INV_X1 _04790_ (.A(_00799_),
    .ZN(\lut.gen_sub_units_scm.__5.sub_unit_i.cg_we_global.en_i ));
 NOR2_X1 _04791_ (.A1(_00665_),
    .A2(_00799_),
    .ZN(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__0.cg_i.en_i ));
 NOR2_X1 _04792_ (.A1(_00668_),
    .A2(_00799_),
    .ZN(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__1.cg_i.en_i ));
 NOR2_X1 _04793_ (.A1(_00671_),
    .A2(_00799_),
    .ZN(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__2.cg_i.en_i ));
 NOR2_X1 _04794_ (.A1(_00673_),
    .A2(_00799_),
    .ZN(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__3.cg_i.en_i ));
 NOR2_X1 _04795_ (.A1(_00678_),
    .A2(_00799_),
    .ZN(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__4.cg_i.en_i ));
 NOR2_X1 _04796_ (.A1(_00680_),
    .A2(_00799_),
    .ZN(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__5.cg_i.en_i ));
 NOR2_X1 _04797_ (.A1(_00681_),
    .A2(_00799_),
    .ZN(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__6.cg_i.en_i ));
 NOR2_X1 _04798_ (.A1(_00682_),
    .A2(_00799_),
    .ZN(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__7.cg_i.en_i ));
 NOR2_X1 _04799_ (.A1(_00686_),
    .A2(_00799_),
    .ZN(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__8.cg_i.en_i ));
 BUF_X4 wire153 (.A(net155),
    .Z(net153));
 NOR2_X1 _04801_ (.A1(_00688_),
    .A2(_00799_),
    .ZN(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__9.cg_i.en_i ));
 NOR2_X1 _04802_ (.A1(_00689_),
    .A2(_00799_),
    .ZN(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__10.cg_i.en_i ));
 NOR2_X1 _04803_ (.A1(_00690_),
    .A2(_00799_),
    .ZN(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__11.cg_i.en_i ));
 NOR2_X1 _04804_ (.A1(_00693_),
    .A2(_00799_),
    .ZN(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__12.cg_i.en_i ));
 NOR2_X1 _04805_ (.A1(_00694_),
    .A2(_00799_),
    .ZN(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__13.cg_i.en_i ));
 NOR2_X1 _04806_ (.A1(_00695_),
    .A2(_00799_),
    .ZN(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__14.cg_i.en_i ));
 NOR2_X1 _04807_ (.A1(_00696_),
    .A2(_00799_),
    .ZN(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__15.cg_i.en_i ));
 NOR2_X1 _04808_ (.A1(_00699_),
    .A2(_00799_),
    .ZN(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__16.cg_i.en_i ));
 NOR2_X1 _04809_ (.A1(_00700_),
    .A2(_00799_),
    .ZN(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__17.cg_i.en_i ));
 NOR2_X1 _04810_ (.A1(_00703_),
    .A2(_00799_),
    .ZN(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__18.cg_i.en_i ));
 BUF_X4 wire152 (.A(_01046_),
    .Z(net152));
 NOR2_X1 _04812_ (.A1(_00707_),
    .A2(_00799_),
    .ZN(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__19.cg_i.en_i ));
 NOR2_X1 _04813_ (.A1(_00709_),
    .A2(_00799_),
    .ZN(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__20.cg_i.en_i ));
 NOR2_X1 _04814_ (.A1(_00711_),
    .A2(_00799_),
    .ZN(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__21.cg_i.en_i ));
 NOR2_X1 _04815_ (.A1(_00712_),
    .A2(_00799_),
    .ZN(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__22.cg_i.en_i ));
 NOR2_X1 _04816_ (.A1(_00713_),
    .A2(_00799_),
    .ZN(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__23.cg_i.en_i ));
 NOR2_X1 _04817_ (.A1(_00714_),
    .A2(_00799_),
    .ZN(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__24.cg_i.en_i ));
 NOR2_X1 _04818_ (.A1(_00715_),
    .A2(_00799_),
    .ZN(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__25.cg_i.en_i ));
 NOR2_X1 _04819_ (.A1(_00716_),
    .A2(_00799_),
    .ZN(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__26.cg_i.en_i ));
 NOR2_X1 _04820_ (.A1(_00717_),
    .A2(_00799_),
    .ZN(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__27.cg_i.en_i ));
 NOR2_X1 _04821_ (.A1(_00718_),
    .A2(_00799_),
    .ZN(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__28.cg_i.en_i ));
 NOR2_X1 _04822_ (.A1(_00719_),
    .A2(_00799_),
    .ZN(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__29.cg_i.en_i ));
 NOR2_X1 _04823_ (.A1(_00720_),
    .A2(_00799_),
    .ZN(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__30.cg_i.en_i ));
 NOR2_X1 _04824_ (.A1(_00721_),
    .A2(_00799_),
    .ZN(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__31.cg_i.en_i ));
 NAND2_X4 _04825_ (.A1(_00765_),
    .A2(_00790_),
    .ZN(_00803_));
 BUF_X4 max_cap151 (.A(_01046_),
    .Z(net151));
 INV_X1 _04827_ (.A(_00803_),
    .ZN(\lut.gen_sub_units_scm.__4.sub_unit_i.cg_we_global.en_i ));
 NOR2_X1 _04828_ (.A1(_00665_),
    .A2(_00803_),
    .ZN(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__0.cg_i.en_i ));
 NOR2_X1 _04829_ (.A1(_00668_),
    .A2(_00803_),
    .ZN(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__1.cg_i.en_i ));
 NOR2_X1 _04830_ (.A1(_00671_),
    .A2(_00803_),
    .ZN(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__2.cg_i.en_i ));
 NOR2_X1 _04831_ (.A1(_00673_),
    .A2(_00803_),
    .ZN(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__3.cg_i.en_i ));
 NOR2_X1 _04832_ (.A1(_00678_),
    .A2(_00803_),
    .ZN(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__4.cg_i.en_i ));
 NOR2_X1 _04833_ (.A1(_00680_),
    .A2(_00803_),
    .ZN(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__5.cg_i.en_i ));
 NOR2_X1 _04834_ (.A1(_00681_),
    .A2(_00803_),
    .ZN(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__6.cg_i.en_i ));
 NOR2_X1 _04835_ (.A1(_00682_),
    .A2(_00803_),
    .ZN(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__7.cg_i.en_i ));
 NOR2_X1 _04836_ (.A1(_00686_),
    .A2(_00803_),
    .ZN(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__8.cg_i.en_i ));
 BUF_X4 max_cap150 (.A(_01046_),
    .Z(net150));
 NOR2_X1 _04838_ (.A1(_00688_),
    .A2(_00803_),
    .ZN(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__9.cg_i.en_i ));
 NOR2_X1 _04839_ (.A1(_00689_),
    .A2(_00803_),
    .ZN(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__10.cg_i.en_i ));
 NOR2_X1 _04840_ (.A1(_00690_),
    .A2(_00803_),
    .ZN(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__11.cg_i.en_i ));
 NOR2_X1 _04841_ (.A1(_00693_),
    .A2(_00803_),
    .ZN(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__12.cg_i.en_i ));
 NOR2_X1 _04842_ (.A1(_00694_),
    .A2(_00803_),
    .ZN(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__13.cg_i.en_i ));
 NOR2_X1 _04843_ (.A1(_00695_),
    .A2(_00803_),
    .ZN(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__14.cg_i.en_i ));
 NOR2_X1 _04844_ (.A1(_00696_),
    .A2(_00803_),
    .ZN(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__15.cg_i.en_i ));
 NOR2_X1 _04845_ (.A1(_00699_),
    .A2(_00803_),
    .ZN(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__16.cg_i.en_i ));
 NOR2_X1 _04846_ (.A1(_00700_),
    .A2(_00803_),
    .ZN(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__17.cg_i.en_i ));
 NOR2_X1 _04847_ (.A1(_00703_),
    .A2(_00803_),
    .ZN(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__18.cg_i.en_i ));
 BUF_X8 max_cap149 (.A(net150),
    .Z(net149));
 NOR2_X1 _04849_ (.A1(_00707_),
    .A2(_00803_),
    .ZN(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__19.cg_i.en_i ));
 NOR2_X1 _04850_ (.A1(_00709_),
    .A2(_00803_),
    .ZN(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__20.cg_i.en_i ));
 NOR2_X1 _04851_ (.A1(_00711_),
    .A2(_00803_),
    .ZN(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__21.cg_i.en_i ));
 NOR2_X1 _04852_ (.A1(_00712_),
    .A2(_00803_),
    .ZN(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__22.cg_i.en_i ));
 NOR2_X1 _04853_ (.A1(_00713_),
    .A2(_00803_),
    .ZN(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__23.cg_i.en_i ));
 NOR2_X1 _04854_ (.A1(_00714_),
    .A2(_00803_),
    .ZN(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__24.cg_i.en_i ));
 NOR2_X1 _04855_ (.A1(_00715_),
    .A2(_00803_),
    .ZN(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__25.cg_i.en_i ));
 NOR2_X1 _04856_ (.A1(_00716_),
    .A2(_00803_),
    .ZN(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__26.cg_i.en_i ));
 NOR2_X1 _04857_ (.A1(_00717_),
    .A2(_00803_),
    .ZN(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__27.cg_i.en_i ));
 NOR2_X1 _04858_ (.A1(_00718_),
    .A2(_00803_),
    .ZN(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__28.cg_i.en_i ));
 NOR2_X1 _04859_ (.A1(_00719_),
    .A2(_00803_),
    .ZN(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__29.cg_i.en_i ));
 NOR2_X1 _04860_ (.A1(_00720_),
    .A2(_00803_),
    .ZN(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__30.cg_i.en_i ));
 NOR2_X1 _04861_ (.A1(_00721_),
    .A2(_00803_),
    .ZN(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__31.cg_i.en_i ));
 NOR3_X4 _04862_ (.A1(net20),
    .A2(net19),
    .A3(_00789_),
    .ZN(_00807_));
 NAND3_X4 _04863_ (.A1(net18),
    .A2(net17),
    .A3(_00807_),
    .ZN(_00808_));
 BUF_X8 max_cap148 (.A(net151),
    .Z(net148));
 INV_X1 _04865_ (.A(_00808_),
    .ZN(\lut.gen_sub_units_scm.__3.sub_unit_i.cg_we_global.en_i ));
 NOR2_X1 _04866_ (.A1(_00665_),
    .A2(_00808_),
    .ZN(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__0.cg_i.en_i ));
 NOR2_X1 _04867_ (.A1(_00668_),
    .A2(_00808_),
    .ZN(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__1.cg_i.en_i ));
 NOR2_X1 _04868_ (.A1(_00671_),
    .A2(_00808_),
    .ZN(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__2.cg_i.en_i ));
 NOR2_X1 _04869_ (.A1(_00673_),
    .A2(_00808_),
    .ZN(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__3.cg_i.en_i ));
 NOR2_X1 _04870_ (.A1(_00678_),
    .A2(_00808_),
    .ZN(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__4.cg_i.en_i ));
 NOR2_X1 _04871_ (.A1(_00680_),
    .A2(_00808_),
    .ZN(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__5.cg_i.en_i ));
 NOR2_X1 _04872_ (.A1(_00681_),
    .A2(_00808_),
    .ZN(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__6.cg_i.en_i ));
 NOR2_X1 _04873_ (.A1(_00682_),
    .A2(_00808_),
    .ZN(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__7.cg_i.en_i ));
 NOR2_X1 _04874_ (.A1(_00686_),
    .A2(_00808_),
    .ZN(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__8.cg_i.en_i ));
 BUF_X4 max_cap147 (.A(net151),
    .Z(net147));
 NOR2_X1 _04876_ (.A1(_00688_),
    .A2(_00808_),
    .ZN(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__9.cg_i.en_i ));
 NOR2_X1 _04877_ (.A1(_00689_),
    .A2(_00808_),
    .ZN(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__10.cg_i.en_i ));
 NOR2_X1 _04878_ (.A1(_00690_),
    .A2(_00808_),
    .ZN(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__11.cg_i.en_i ));
 NOR2_X1 _04879_ (.A1(_00693_),
    .A2(_00808_),
    .ZN(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__12.cg_i.en_i ));
 NOR2_X1 _04880_ (.A1(_00694_),
    .A2(_00808_),
    .ZN(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__13.cg_i.en_i ));
 NOR2_X1 _04881_ (.A1(_00695_),
    .A2(_00808_),
    .ZN(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__14.cg_i.en_i ));
 NOR2_X1 _04882_ (.A1(_00696_),
    .A2(_00808_),
    .ZN(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__15.cg_i.en_i ));
 NOR2_X1 _04883_ (.A1(_00699_),
    .A2(_00808_),
    .ZN(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__16.cg_i.en_i ));
 NOR2_X1 _04884_ (.A1(_00700_),
    .A2(_00808_),
    .ZN(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__17.cg_i.en_i ));
 NOR2_X1 _04885_ (.A1(_00703_),
    .A2(_00808_),
    .ZN(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__18.cg_i.en_i ));
 BUF_X8 max_cap146 (.A(_01050_),
    .Z(net146));
 NOR2_X1 _04887_ (.A1(_00707_),
    .A2(_00808_),
    .ZN(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__19.cg_i.en_i ));
 NOR2_X1 _04888_ (.A1(_00709_),
    .A2(_00808_),
    .ZN(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__20.cg_i.en_i ));
 NOR2_X1 _04889_ (.A1(_00711_),
    .A2(_00808_),
    .ZN(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__21.cg_i.en_i ));
 NOR2_X1 _04890_ (.A1(_00712_),
    .A2(_00808_),
    .ZN(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__22.cg_i.en_i ));
 NOR2_X1 _04891_ (.A1(_00713_),
    .A2(_00808_),
    .ZN(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__23.cg_i.en_i ));
 NOR2_X1 _04892_ (.A1(_00714_),
    .A2(_00808_),
    .ZN(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__24.cg_i.en_i ));
 NOR2_X1 _04893_ (.A1(_00715_),
    .A2(_00808_),
    .ZN(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__25.cg_i.en_i ));
 NOR2_X1 _04894_ (.A1(_00716_),
    .A2(_00808_),
    .ZN(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__26.cg_i.en_i ));
 NOR2_X1 _04895_ (.A1(_00717_),
    .A2(_00808_),
    .ZN(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__27.cg_i.en_i ));
 NOR2_X1 _04896_ (.A1(_00718_),
    .A2(_00808_),
    .ZN(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__28.cg_i.en_i ));
 NOR2_X1 _04897_ (.A1(_00719_),
    .A2(_00808_),
    .ZN(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__29.cg_i.en_i ));
 NOR2_X1 _04898_ (.A1(_00720_),
    .A2(_00808_),
    .ZN(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__30.cg_i.en_i ));
 NOR2_X1 _04899_ (.A1(_00721_),
    .A2(_00808_),
    .ZN(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__31.cg_i.en_i ));
 NAND2_X4 _04900_ (.A1(_00723_),
    .A2(_00807_),
    .ZN(_00812_));
 BUF_X8 max_cap145 (.A(_01050_),
    .Z(net145));
 INV_X1 _04902_ (.A(_00812_),
    .ZN(\lut.gen_sub_units_scm.__2.sub_unit_i.cg_we_global.en_i ));
 NOR2_X1 _04903_ (.A1(_00665_),
    .A2(_00812_),
    .ZN(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__0.cg_i.en_i ));
 NOR2_X1 _04904_ (.A1(_00668_),
    .A2(_00812_),
    .ZN(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__1.cg_i.en_i ));
 NOR2_X1 _04905_ (.A1(_00671_),
    .A2(_00812_),
    .ZN(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__2.cg_i.en_i ));
 NOR2_X1 _04906_ (.A1(_00673_),
    .A2(_00812_),
    .ZN(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__3.cg_i.en_i ));
 NOR2_X1 _04907_ (.A1(_00678_),
    .A2(_00812_),
    .ZN(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__4.cg_i.en_i ));
 NOR2_X1 _04908_ (.A1(_00680_),
    .A2(_00812_),
    .ZN(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__5.cg_i.en_i ));
 NOR2_X1 _04909_ (.A1(_00681_),
    .A2(_00812_),
    .ZN(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__6.cg_i.en_i ));
 NOR2_X1 _04910_ (.A1(_00682_),
    .A2(_00812_),
    .ZN(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__7.cg_i.en_i ));
 NOR2_X1 _04911_ (.A1(_00686_),
    .A2(_00812_),
    .ZN(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__8.cg_i.en_i ));
 BUF_X8 max_cap144 (.A(net145),
    .Z(net144));
 NOR2_X1 _04913_ (.A1(_00688_),
    .A2(_00812_),
    .ZN(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__9.cg_i.en_i ));
 NOR2_X1 _04914_ (.A1(_00689_),
    .A2(_00812_),
    .ZN(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__10.cg_i.en_i ));
 NOR2_X1 _04915_ (.A1(_00690_),
    .A2(_00812_),
    .ZN(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__11.cg_i.en_i ));
 NOR2_X1 _04916_ (.A1(_00693_),
    .A2(_00812_),
    .ZN(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__12.cg_i.en_i ));
 NOR2_X1 _04917_ (.A1(_00694_),
    .A2(_00812_),
    .ZN(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__13.cg_i.en_i ));
 NOR2_X1 _04918_ (.A1(_00695_),
    .A2(_00812_),
    .ZN(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__14.cg_i.en_i ));
 NOR2_X1 _04919_ (.A1(_00696_),
    .A2(_00812_),
    .ZN(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__15.cg_i.en_i ));
 NOR2_X1 _04920_ (.A1(_00699_),
    .A2(_00812_),
    .ZN(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__16.cg_i.en_i ));
 NOR2_X1 _04921_ (.A1(_00700_),
    .A2(_00812_),
    .ZN(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__17.cg_i.en_i ));
 NOR2_X1 _04922_ (.A1(_00703_),
    .A2(_00812_),
    .ZN(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__18.cg_i.en_i ));
 BUF_X8 max_cap143 (.A(net145),
    .Z(net143));
 NOR2_X1 _04924_ (.A1(_00707_),
    .A2(_00812_),
    .ZN(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__19.cg_i.en_i ));
 NOR2_X1 _04925_ (.A1(_00709_),
    .A2(_00812_),
    .ZN(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__20.cg_i.en_i ));
 NOR2_X1 _04926_ (.A1(_00711_),
    .A2(_00812_),
    .ZN(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__21.cg_i.en_i ));
 NOR2_X1 _04927_ (.A1(_00712_),
    .A2(_00812_),
    .ZN(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__22.cg_i.en_i ));
 NOR2_X1 _04928_ (.A1(_00713_),
    .A2(_00812_),
    .ZN(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__23.cg_i.en_i ));
 NOR2_X1 _04929_ (.A1(_00714_),
    .A2(_00812_),
    .ZN(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__24.cg_i.en_i ));
 NOR2_X1 _04930_ (.A1(_00715_),
    .A2(_00812_),
    .ZN(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__25.cg_i.en_i ));
 NOR2_X1 _04931_ (.A1(_00716_),
    .A2(_00812_),
    .ZN(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__26.cg_i.en_i ));
 NOR2_X1 _04932_ (.A1(_00717_),
    .A2(_00812_),
    .ZN(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__27.cg_i.en_i ));
 NOR2_X1 _04933_ (.A1(_00718_),
    .A2(_00812_),
    .ZN(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__28.cg_i.en_i ));
 NOR2_X1 _04934_ (.A1(_00719_),
    .A2(_00812_),
    .ZN(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__29.cg_i.en_i ));
 NOR2_X1 _04935_ (.A1(_00720_),
    .A2(_00812_),
    .ZN(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__30.cg_i.en_i ));
 NOR2_X1 _04936_ (.A1(_00721_),
    .A2(_00812_),
    .ZN(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__31.cg_i.en_i ));
 NAND2_X4 _04937_ (.A1(_00760_),
    .A2(_00807_),
    .ZN(_00816_));
 BUF_X8 max_cap142 (.A(net145),
    .Z(net142));
 INV_X1 _04939_ (.A(_00816_),
    .ZN(\lut.gen_sub_units_scm.__1.sub_unit_i.cg_we_global.en_i ));
 NOR2_X1 _04940_ (.A1(_00665_),
    .A2(_00816_),
    .ZN(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__0.cg_i.en_i ));
 NOR2_X1 _04941_ (.A1(_00668_),
    .A2(_00816_),
    .ZN(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__1.cg_i.en_i ));
 NOR2_X1 _04942_ (.A1(_00671_),
    .A2(_00816_),
    .ZN(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__2.cg_i.en_i ));
 NOR2_X1 _04943_ (.A1(_00673_),
    .A2(_00816_),
    .ZN(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__3.cg_i.en_i ));
 NOR2_X1 _04944_ (.A1(_00678_),
    .A2(_00816_),
    .ZN(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__4.cg_i.en_i ));
 NOR2_X1 _04945_ (.A1(_00680_),
    .A2(_00816_),
    .ZN(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__5.cg_i.en_i ));
 NOR2_X1 _04946_ (.A1(_00681_),
    .A2(_00816_),
    .ZN(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__6.cg_i.en_i ));
 NOR2_X1 _04947_ (.A1(_00682_),
    .A2(_00816_),
    .ZN(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__7.cg_i.en_i ));
 NOR2_X1 _04948_ (.A1(_00686_),
    .A2(_00816_),
    .ZN(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__8.cg_i.en_i ));
 BUF_X8 wire141 (.A(_01050_),
    .Z(net141));
 NOR2_X1 _04950_ (.A1(_00688_),
    .A2(_00816_),
    .ZN(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__9.cg_i.en_i ));
 NOR2_X1 _04951_ (.A1(_00689_),
    .A2(_00816_),
    .ZN(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__10.cg_i.en_i ));
 NOR2_X1 _04952_ (.A1(_00690_),
    .A2(_00816_),
    .ZN(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__11.cg_i.en_i ));
 NOR2_X1 _04953_ (.A1(_00693_),
    .A2(_00816_),
    .ZN(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__12.cg_i.en_i ));
 NOR2_X1 _04954_ (.A1(_00694_),
    .A2(_00816_),
    .ZN(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__13.cg_i.en_i ));
 NOR2_X1 _04955_ (.A1(_00695_),
    .A2(_00816_),
    .ZN(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__14.cg_i.en_i ));
 NOR2_X1 _04956_ (.A1(_00696_),
    .A2(_00816_),
    .ZN(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__15.cg_i.en_i ));
 NOR2_X1 _04957_ (.A1(_00699_),
    .A2(_00816_),
    .ZN(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__16.cg_i.en_i ));
 NOR2_X1 _04958_ (.A1(_00700_),
    .A2(_00816_),
    .ZN(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__17.cg_i.en_i ));
 NOR2_X1 _04959_ (.A1(_00703_),
    .A2(_00816_),
    .ZN(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__18.cg_i.en_i ));
 BUF_X8 max_cap140 (.A(net146),
    .Z(net140));
 NOR2_X1 _04961_ (.A1(_00707_),
    .A2(_00816_),
    .ZN(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__19.cg_i.en_i ));
 NOR2_X1 _04962_ (.A1(_00709_),
    .A2(_00816_),
    .ZN(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__20.cg_i.en_i ));
 NOR2_X1 _04963_ (.A1(_00711_),
    .A2(_00816_),
    .ZN(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__21.cg_i.en_i ));
 NOR2_X1 _04964_ (.A1(_00712_),
    .A2(_00816_),
    .ZN(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__22.cg_i.en_i ));
 NOR2_X1 _04965_ (.A1(_00713_),
    .A2(_00816_),
    .ZN(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__23.cg_i.en_i ));
 NOR2_X1 _04966_ (.A1(_00714_),
    .A2(_00816_),
    .ZN(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__24.cg_i.en_i ));
 NOR2_X1 _04967_ (.A1(_00715_),
    .A2(_00816_),
    .ZN(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__25.cg_i.en_i ));
 NOR2_X1 _04968_ (.A1(_00716_),
    .A2(_00816_),
    .ZN(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__26.cg_i.en_i ));
 NOR2_X1 _04969_ (.A1(_00717_),
    .A2(_00816_),
    .ZN(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__27.cg_i.en_i ));
 NOR2_X1 _04970_ (.A1(_00718_),
    .A2(_00816_),
    .ZN(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__28.cg_i.en_i ));
 NOR2_X1 _04971_ (.A1(_00719_),
    .A2(_00816_),
    .ZN(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__29.cg_i.en_i ));
 NOR2_X1 _04972_ (.A1(_00720_),
    .A2(_00816_),
    .ZN(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__30.cg_i.en_i ));
 NOR2_X1 _04973_ (.A1(_00721_),
    .A2(_00816_),
    .ZN(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__31.cg_i.en_i ));
 NAND2_X4 _04974_ (.A1(_00765_),
    .A2(_00807_),
    .ZN(_00820_));
 BUF_X4 max_cap139 (.A(_01057_),
    .Z(net139));
 INV_X1 _04976_ (.A(_00820_),
    .ZN(\lut.gen_sub_units_scm.__0.sub_unit_i.cg_we_global.en_i ));
 NOR2_X1 _04977_ (.A1(_00665_),
    .A2(_00820_),
    .ZN(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__0.cg_i.en_i ));
 NOR2_X1 _04978_ (.A1(_00668_),
    .A2(_00820_),
    .ZN(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__1.cg_i.en_i ));
 NOR2_X1 _04979_ (.A1(_00671_),
    .A2(_00820_),
    .ZN(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__2.cg_i.en_i ));
 NOR2_X1 _04980_ (.A1(_00673_),
    .A2(_00820_),
    .ZN(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__3.cg_i.en_i ));
 NOR2_X1 _04981_ (.A1(_00678_),
    .A2(_00820_),
    .ZN(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__4.cg_i.en_i ));
 NOR2_X1 _04982_ (.A1(_00680_),
    .A2(_00820_),
    .ZN(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__5.cg_i.en_i ));
 NOR2_X1 _04983_ (.A1(_00681_),
    .A2(_00820_),
    .ZN(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__6.cg_i.en_i ));
 NOR2_X1 _04984_ (.A1(_00682_),
    .A2(_00820_),
    .ZN(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__7.cg_i.en_i ));
 NOR2_X1 _04985_ (.A1(_00686_),
    .A2(_00820_),
    .ZN(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__8.cg_i.en_i ));
 BUF_X8 max_cap138 (.A(net139),
    .Z(net138));
 NOR2_X1 _04987_ (.A1(_00688_),
    .A2(_00820_),
    .ZN(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__9.cg_i.en_i ));
 NOR2_X1 _04988_ (.A1(_00689_),
    .A2(_00820_),
    .ZN(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__10.cg_i.en_i ));
 NOR2_X1 _04989_ (.A1(_00690_),
    .A2(_00820_),
    .ZN(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__11.cg_i.en_i ));
 NOR2_X1 _04990_ (.A1(_00693_),
    .A2(_00820_),
    .ZN(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__12.cg_i.en_i ));
 NOR2_X1 _04991_ (.A1(_00694_),
    .A2(_00820_),
    .ZN(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__13.cg_i.en_i ));
 NOR2_X1 _04992_ (.A1(_00695_),
    .A2(_00820_),
    .ZN(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__14.cg_i.en_i ));
 NOR2_X1 _04993_ (.A1(_00696_),
    .A2(_00820_),
    .ZN(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__15.cg_i.en_i ));
 NOR2_X1 _04994_ (.A1(_00699_),
    .A2(_00820_),
    .ZN(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__16.cg_i.en_i ));
 NOR2_X1 _04995_ (.A1(_00700_),
    .A2(_00820_),
    .ZN(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__17.cg_i.en_i ));
 NOR2_X1 _04996_ (.A1(_00703_),
    .A2(_00820_),
    .ZN(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__18.cg_i.en_i ));
 BUF_X4 max_cap137 (.A(net138),
    .Z(net137));
 NOR2_X1 _04998_ (.A1(_00707_),
    .A2(_00820_),
    .ZN(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__19.cg_i.en_i ));
 NOR2_X1 _04999_ (.A1(_00709_),
    .A2(_00820_),
    .ZN(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__20.cg_i.en_i ));
 NOR2_X1 _05000_ (.A1(_00711_),
    .A2(_00820_),
    .ZN(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__21.cg_i.en_i ));
 NOR2_X1 _05001_ (.A1(_00712_),
    .A2(_00820_),
    .ZN(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__22.cg_i.en_i ));
 NOR2_X1 _05002_ (.A1(_00713_),
    .A2(_00820_),
    .ZN(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__23.cg_i.en_i ));
 NOR2_X1 _05003_ (.A1(_00714_),
    .A2(_00820_),
    .ZN(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__24.cg_i.en_i ));
 NOR2_X1 _05004_ (.A1(_00715_),
    .A2(_00820_),
    .ZN(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__25.cg_i.en_i ));
 NOR2_X1 _05005_ (.A1(_00716_),
    .A2(_00820_),
    .ZN(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__26.cg_i.en_i ));
 NOR2_X1 _05006_ (.A1(_00717_),
    .A2(_00820_),
    .ZN(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__27.cg_i.en_i ));
 NOR2_X1 _05007_ (.A1(_00718_),
    .A2(_00820_),
    .ZN(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__28.cg_i.en_i ));
 NOR2_X1 _05008_ (.A1(_00719_),
    .A2(_00820_),
    .ZN(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__29.cg_i.en_i ));
 NOR2_X1 _05009_ (.A1(_00720_),
    .A2(_00820_),
    .ZN(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__30.cg_i.en_i ));
 NOR2_X1 _05010_ (.A1(_00721_),
    .A2(_00820_),
    .ZN(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__31.cg_i.en_i ));
 BUF_X4 max_cap136 (.A(net138),
    .Z(net136));
 INV_X1 _05012_ (.A(\caddr_q[4] ),
    .ZN(_00825_));
 NAND4_X1 _05013_ (.A1(\caddr_q[1] ),
    .A2(\caddr_q[0] ),
    .A3(\caddr_q[3] ),
    .A4(\caddr_q[2] ),
    .ZN(_00826_));
 OR2_X4 _05014_ (.A1(_00825_),
    .A2(_00826_),
    .ZN(_00827_));
 BUF_X4 wire135 (.A(_01057_),
    .Z(net135));
 BUF_X4 max_cap134 (.A(_01057_),
    .Z(net134));
 AND2_X1 _05017_ (.A1(net6),
    .A2(_00827_),
    .ZN(_00830_));
 AND2_X1 _05018_ (.A1(_04253_),
    .A2(_00830_),
    .ZN(\result_int_n[0] ));
 NAND2_X4 _05019_ (.A1(net6),
    .A2(_00827_),
    .ZN(_00831_));
 BUF_X4 max_cap133 (.A(_01057_),
    .Z(net133));
 NOR2_X1 _05021_ (.A1(_04198_),
    .A2(_00831_),
    .ZN(\result_int_n[1] ));
 AND2_X1 _05022_ (.A1(_04200_),
    .A2(_00830_),
    .ZN(\result_int_n[2] ));
 BUF_X8 max_cap132 (.A(net134),
    .Z(net132));
 XNOR2_X1 _05024_ (.A(_04257_),
    .B(_04199_),
    .ZN(_00834_));
 NOR2_X1 _05025_ (.A1(_00831_),
    .A2(_00834_),
    .ZN(\result_int_n[3] ));
 INV_X1 _05026_ (.A(_04256_),
    .ZN(_00835_));
 AOI21_X1 _05027_ (.A(_04254_),
    .B1(_04255_),
    .B2(_04197_),
    .ZN(_00836_));
 INV_X1 _05028_ (.A(_04257_),
    .ZN(_00837_));
 OAI21_X1 _05029_ (.A(_00835_),
    .B1(_00836_),
    .B2(_00837_),
    .ZN(_04201_));
 AND2_X1 _05030_ (.A1(_04203_),
    .A2(_00830_),
    .ZN(\result_int_n[4] ));
 XNOR2_X1 _05031_ (.A(_04261_),
    .B(_04202_),
    .ZN(_00838_));
 NOR2_X1 _05032_ (.A1(_00831_),
    .A2(_00838_),
    .ZN(\result_int_n[5] ));
 NAND2_X1 _05033_ (.A1(_04261_),
    .A2(_04259_),
    .ZN(_00839_));
 NOR3_X1 _05034_ (.A1(_00837_),
    .A2(_00836_),
    .A3(_00839_),
    .ZN(_00840_));
 INV_X1 _05035_ (.A(_04261_),
    .ZN(_00841_));
 AOI21_X1 _05036_ (.A(_04258_),
    .B1(_04259_),
    .B2(_04256_),
    .ZN(_00842_));
 NOR2_X1 _05037_ (.A1(_00841_),
    .A2(_00842_),
    .ZN(_00843_));
 NOR3_X2 _05038_ (.A1(_04260_),
    .A2(_00840_),
    .A3(_00843_),
    .ZN(_04204_));
 NOR2_X1 _05039_ (.A1(_04208_),
    .A2(_00831_),
    .ZN(\result_int_n[6] ));
 XOR2_X1 _05040_ (.A(_04207_),
    .B(_04265_),
    .Z(_00844_));
 NOR2_X1 _05041_ (.A1(_00831_),
    .A2(_00844_),
    .ZN(\result_int_n[7] ));
 AOI21_X1 _05042_ (.A(_04264_),
    .B1(_04262_),
    .B2(_04265_),
    .ZN(_00845_));
 NAND2_X1 _05043_ (.A1(_04265_),
    .A2(_04263_),
    .ZN(_00846_));
 OAI21_X1 _05044_ (.A(_00845_),
    .B1(_00846_),
    .B2(_04204_),
    .ZN(_04209_));
 AND2_X1 _05045_ (.A1(_04211_),
    .A2(_00830_),
    .ZN(\result_int_n[8] ));
 BUF_X8 max_cap131 (.A(net134),
    .Z(net131));
 XNOR2_X1 _05047_ (.A(_04269_),
    .B(_04210_),
    .ZN(_00848_));
 NOR2_X1 _05048_ (.A1(_00831_),
    .A2(_00848_),
    .ZN(\result_int_n[9] ));
 AOI21_X1 _05049_ (.A(_04266_),
    .B1(_04209_),
    .B2(_04267_),
    .ZN(_00849_));
 INV_X1 _05050_ (.A(_00849_),
    .ZN(_00850_));
 AOI21_X1 _05051_ (.A(_04268_),
    .B1(_00850_),
    .B2(_04269_),
    .ZN(_04212_));
 NOR2_X1 _05052_ (.A1(_04216_),
    .A2(_00831_),
    .ZN(\result_int_n[10] ));
 BUF_X32 max_cap130 (.A(_01064_),
    .Z(net130));
 XOR2_X1 _05054_ (.A(_04215_),
    .B(_04273_),
    .Z(_00852_));
 NOR2_X1 _05055_ (.A1(_00831_),
    .A2(_00852_),
    .ZN(\result_int_n[11] ));
 AOI21_X1 _05056_ (.A(_04268_),
    .B1(_04266_),
    .B2(_04269_),
    .ZN(_00853_));
 NAND2_X1 _05057_ (.A1(_04273_),
    .A2(_04271_),
    .ZN(_00854_));
 NOR2_X1 _05058_ (.A1(_00853_),
    .A2(_00854_),
    .ZN(_00855_));
 AOI21_X1 _05059_ (.A(_04272_),
    .B1(_04270_),
    .B2(_04273_),
    .ZN(_00856_));
 NAND4_X1 _05060_ (.A1(_04269_),
    .A2(_04273_),
    .A3(_04267_),
    .A4(_04271_),
    .ZN(_00857_));
 OAI21_X1 _05061_ (.A(_00856_),
    .B1(_00857_),
    .B2(_00845_),
    .ZN(_00858_));
 NOR2_X1 _05062_ (.A1(_00855_),
    .A2(_00858_),
    .ZN(_00859_));
 OR2_X1 _05063_ (.A1(_00846_),
    .A2(_00857_),
    .ZN(_00860_));
 OAI21_X2 _05064_ (.A(_00859_),
    .B1(_00860_),
    .B2(_04204_),
    .ZN(_00861_));
 INV_X1 _05065_ (.A(_00861_),
    .ZN(_04217_));
 NOR2_X1 _05066_ (.A1(_04220_),
    .A2(_00831_),
    .ZN(\result_int_n[12] ));
 XOR2_X1 _05067_ (.A(_04219_),
    .B(_04277_),
    .Z(_00862_));
 NOR2_X1 _05068_ (.A1(_00831_),
    .A2(_00862_),
    .ZN(\result_int_n[13] ));
 AOI21_X1 _05069_ (.A(_04276_),
    .B1(_04274_),
    .B2(_04277_),
    .ZN(_00863_));
 NAND3_X1 _05070_ (.A1(_04277_),
    .A2(_04275_),
    .A3(_00861_),
    .ZN(_00864_));
 AND2_X1 _05071_ (.A1(_00863_),
    .A2(_00864_),
    .ZN(_04221_));
 NOR2_X1 _05072_ (.A1(_04224_),
    .A2(_00831_),
    .ZN(\result_int_n[14] ));
 XOR2_X1 _05073_ (.A(_04223_),
    .B(_04281_),
    .Z(_00865_));
 NOR2_X1 _05074_ (.A1(_00831_),
    .A2(_00865_),
    .ZN(\result_int_n[15] ));
 AND4_X1 _05075_ (.A1(_04277_),
    .A2(_04281_),
    .A3(_04275_),
    .A4(_04279_),
    .ZN(_00866_));
 INV_X1 _05076_ (.A(_04278_),
    .ZN(_00867_));
 INV_X1 _05077_ (.A(_04279_),
    .ZN(_00868_));
 OAI21_X1 _05078_ (.A(_00867_),
    .B1(_00863_),
    .B2(_00868_),
    .ZN(_00869_));
 AOI221_X2 _05079_ (.A(_04280_),
    .B1(_00861_),
    .B2(_00866_),
    .C1(_00869_),
    .C2(_04281_),
    .ZN(_00870_));
 INV_X1 _05080_ (.A(_00870_),
    .ZN(_04225_));
 AND2_X1 _05081_ (.A1(_04227_),
    .A2(_00830_),
    .ZN(\result_int_n[16] ));
 XNOR2_X1 _05082_ (.A(_04285_),
    .B(_04226_),
    .ZN(_00871_));
 NOR2_X1 _05083_ (.A1(_00831_),
    .A2(_00871_),
    .ZN(\result_int_n[17] ));
 AND2_X1 _05084_ (.A1(_04285_),
    .A2(_04283_),
    .ZN(_00872_));
 AOI221_X2 _05085_ (.A(_04284_),
    .B1(_04225_),
    .B2(_00872_),
    .C1(_04282_),
    .C2(_04285_),
    .ZN(_04228_));
 NOR2_X1 _05086_ (.A1(_04231_),
    .A2(_00831_),
    .ZN(\result_int_n[18] ));
 XOR2_X1 _05087_ (.A(_04230_),
    .B(_04289_),
    .Z(_00873_));
 NOR2_X1 _05088_ (.A1(_00831_),
    .A2(_00873_),
    .ZN(\result_int_n[19] ));
 INV_X1 _05089_ (.A(_04286_),
    .ZN(_00874_));
 AOI21_X1 _05090_ (.A(_04284_),
    .B1(_04282_),
    .B2(_04285_),
    .ZN(_00875_));
 INV_X1 _05091_ (.A(_04287_),
    .ZN(_00876_));
 OAI21_X1 _05092_ (.A(_00874_),
    .B1(_00875_),
    .B2(_00876_),
    .ZN(_00877_));
 AOI21_X1 _05093_ (.A(_04288_),
    .B1(_00877_),
    .B2(_04289_),
    .ZN(_00878_));
 NAND3_X1 _05094_ (.A1(_04289_),
    .A2(_04287_),
    .A3(_00872_),
    .ZN(_00879_));
 OR2_X1 _05095_ (.A1(_00870_),
    .A2(_00879_),
    .ZN(_00880_));
 AND2_X1 _05096_ (.A1(_00878_),
    .A2(_00880_),
    .ZN(_04232_));
 NOR2_X1 _05097_ (.A1(_04235_),
    .A2(_00831_),
    .ZN(\result_int_n[20] ));
 BUF_X8 max_cap129 (.A(_01081_),
    .Z(net129));
 XOR2_X1 _05099_ (.A(_04234_),
    .B(_04293_),
    .Z(_00882_));
 NOR2_X1 _05100_ (.A1(_00831_),
    .A2(_00882_),
    .ZN(\result_int_n[21] ));
 NOR2_X1 _05101_ (.A1(_04238_),
    .A2(_00831_),
    .ZN(\result_int_n[22] ));
 XNOR2_X1 _05102_ (.A(_04237_),
    .B(_04297_),
    .ZN(_00883_));
 NOR2_X1 _05103_ (.A1(_00831_),
    .A2(_00883_),
    .ZN(\result_int_n[23] ));
 AND2_X1 _05104_ (.A1(_04242_),
    .A2(_00830_),
    .ZN(\result_int_n[24] ));
 XOR2_X1 _05105_ (.A(_04241_),
    .B(_04301_),
    .Z(_00884_));
 NOR2_X1 _05106_ (.A1(_00831_),
    .A2(_00884_),
    .ZN(\result_int_n[25] ));
 NOR2_X1 _05107_ (.A1(_04245_),
    .A2(_00831_),
    .ZN(\result_int_n[26] ));
 XNOR2_X1 _05108_ (.A(_04244_),
    .B(_04305_),
    .ZN(_00885_));
 NOR2_X1 _05109_ (.A1(_00831_),
    .A2(_00885_),
    .ZN(\result_int_n[27] ));
 NOR2_X1 _05110_ (.A1(_04248_),
    .A2(_00831_),
    .ZN(\result_int_n[28] ));
 XNOR2_X1 _05111_ (.A(_04247_),
    .B(_04309_),
    .ZN(_00886_));
 NOR2_X1 _05112_ (.A1(_00831_),
    .A2(_00886_),
    .ZN(\result_int_n[29] ));
 AOI21_X1 _05113_ (.A(_04304_),
    .B1(_04302_),
    .B2(_04305_),
    .ZN(_00887_));
 NAND2_X1 _05114_ (.A1(_04303_),
    .A2(_04305_),
    .ZN(_00888_));
 INV_X1 _05115_ (.A(_04294_),
    .ZN(_00889_));
 AOI21_X1 _05116_ (.A(_04292_),
    .B1(_04290_),
    .B2(_04293_),
    .ZN(_00890_));
 INV_X1 _05117_ (.A(_04295_),
    .ZN(_00891_));
 OAI21_X1 _05118_ (.A(_00889_),
    .B1(_00890_),
    .B2(_00891_),
    .ZN(_00892_));
 AOI21_X1 _05119_ (.A(_04296_),
    .B1(_04297_),
    .B2(_00892_),
    .ZN(_00893_));
 NAND4_X1 _05120_ (.A1(_04293_),
    .A2(_04291_),
    .A3(_04295_),
    .A4(_04297_),
    .ZN(_00894_));
 OAI21_X1 _05121_ (.A(_00893_),
    .B1(_00894_),
    .B2(_00878_),
    .ZN(_00895_));
 NOR3_X1 _05122_ (.A1(_04300_),
    .A2(_04298_),
    .A3(_00895_),
    .ZN(_00896_));
 OR2_X1 _05123_ (.A1(_00879_),
    .A2(_00894_),
    .ZN(_00897_));
 OAI21_X1 _05124_ (.A(_00896_),
    .B1(_00897_),
    .B2(_00870_),
    .ZN(_00898_));
 NOR2_X1 _05125_ (.A1(_04300_),
    .A2(_04301_),
    .ZN(_00899_));
 NOR2_X1 _05126_ (.A1(_04300_),
    .A2(_04299_),
    .ZN(_00900_));
 INV_X1 _05127_ (.A(_04298_),
    .ZN(_00901_));
 AOI21_X1 _05128_ (.A(_00899_),
    .B1(_00900_),
    .B2(_00901_),
    .ZN(_00902_));
 NAND2_X1 _05129_ (.A1(_00898_),
    .A2(_00902_),
    .ZN(_00903_));
 OAI21_X2 _05130_ (.A(_00887_),
    .B1(_00888_),
    .B2(_00903_),
    .ZN(_04246_));
 AND2_X1 _05131_ (.A1(_04307_),
    .A2(_04309_),
    .ZN(_00904_));
 AOI221_X2 _05132_ (.A(_04308_),
    .B1(_04246_),
    .B2(_00904_),
    .C1(_04306_),
    .C2(_04309_),
    .ZN(_04249_));
 NOR2_X1 _05133_ (.A1(_04252_),
    .A2(_00831_),
    .ZN(\result_int_n[30] ));
 XNOR2_X1 _05134_ (.A(\genblk1.gen_int_accumulation.int_adder.int_short_converted[10] ),
    .B(_04251_),
    .ZN(_00905_));
 XNOR2_X1 _05135_ (.A(\genblk1.gen_int_accumulation.int_adder.int_long_i[31] ),
    .B(_00905_),
    .ZN(_00906_));
 NOR2_X1 _05136_ (.A1(_00831_),
    .A2(_00906_),
    .ZN(\result_int_n[31] ));
 INV_X8 _05137_ (.A(net6),
    .ZN(_00907_));
 BUF_X16 max_cap128 (.A(net129),
    .Z(net128));
 BUF_X8 max_cap127 (.A(net129),
    .Z(net127));
 BUF_X8 max_cap126 (.A(_01081_),
    .Z(net126));
 INV_X8 _05141_ (.A(net1),
    .ZN(_00911_));
 BUF_X8 wire125 (.A(_01081_),
    .Z(net125));
 NOR2_X1 _05143_ (.A1(_00907_),
    .A2(_00911_),
    .ZN(\caddr_n[0] ));
 BUF_X8 max_cap124 (.A(net125),
    .Z(net124));
 INV_X2 _05145_ (.A(net2),
    .ZN(_00914_));
 NOR2_X1 _05146_ (.A1(_00907_),
    .A2(_00914_),
    .ZN(\caddr_n[1] ));
 BUF_X8 max_cap123 (.A(net126),
    .Z(net123));
 INV_X2 _05148_ (.A(net3),
    .ZN(_00916_));
 NOR2_X1 _05149_ (.A1(_00907_),
    .A2(_00916_),
    .ZN(\caddr_n[2] ));
 BUF_X8 max_cap122 (.A(_01097_),
    .Z(net122));
 INV_X2 _05151_ (.A(net4),
    .ZN(_00918_));
 NOR2_X1 _05152_ (.A1(_00907_),
    .A2(_00918_),
    .ZN(\caddr_n[3] ));
 BUF_X8 max_cap121 (.A(net122),
    .Z(net121));
 INV_X2 _05154_ (.A(net5),
    .ZN(_00920_));
 NOR2_X1 _05155_ (.A1(_00907_),
    .A2(_00920_),
    .ZN(\caddr_n[4] ));
 NAND2_X4 _05156_ (.A1(net2),
    .A2(_00916_),
    .ZN(_00921_));
 NAND2_X4 _05157_ (.A1(_00918_),
    .A2(net5),
    .ZN(_00922_));
 NOR2_X4 _05158_ (.A1(_00921_),
    .A2(_00922_),
    .ZN(_00923_));
 INV_X1 _05159_ (.A(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[31][0] ),
    .ZN(_00924_));
 BUF_X8 max_cap120 (.A(_01097_),
    .Z(net120));
 AND2_X4 _05161_ (.A1(net1),
    .A2(net8),
    .ZN(_00926_));
 BUF_X8 max_cap119 (.A(_01097_),
    .Z(net119));
 BUF_X8 max_cap118 (.A(_01097_),
    .Z(net118));
 BUF_X8 max_cap117 (.A(net120),
    .Z(net117));
 BUF_X8 max_cap116 (.A(net117),
    .Z(net116));
 BUF_X16 max_cap115 (.A(_01119_),
    .Z(net115));
 BUF_X16 max_cap114 (.A(_01119_),
    .Z(net114));
 AND3_X4 _05168_ (.A1(net7),
    .A2(net10),
    .A3(net9),
    .ZN(_00933_));
 NAND2_X4 _05169_ (.A1(_00926_),
    .A2(_00933_),
    .ZN(_00934_));
 BUF_X16 max_length113 (.A(net114),
    .Z(net113));
 BUF_X8 max_cap112 (.A(_01123_),
    .Z(net112));
 NOR2_X4 _05172_ (.A1(net7),
    .A2(net10),
    .ZN(_00937_));
 BUF_X8 max_cap111 (.A(net112),
    .Z(net111));
 NOR2_X4 _05174_ (.A1(net1),
    .A2(net8),
    .ZN(_00939_));
 BUF_X8 max_cap110 (.A(net111),
    .Z(net110));
 NAND3_X4 _05176_ (.A1(net9),
    .A2(_00937_),
    .A3(_00939_),
    .ZN(_00941_));
 INV_X1 _05177_ (.A(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[4][0] ),
    .ZN(_00942_));
 OAI22_X1 _05178_ (.A1(_00924_),
    .A2(_00934_),
    .B1(_00941_),
    .B2(_00942_),
    .ZN(_00943_));
 INV_X8 _05179_ (.A(net10),
    .ZN(_00944_));
 BUF_X8 max_cap109 (.A(_01123_),
    .Z(net109));
 INV_X16 _05181_ (.A(net9),
    .ZN(_00946_));
 BUF_X8 max_cap108 (.A(_01123_),
    .Z(net108));
 OR2_X4 _05183_ (.A1(net1),
    .A2(net8),
    .ZN(_00948_));
 BUF_X8 max_cap107 (.A(net108),
    .Z(net107));
 NOR4_X4 _05185_ (.A1(net7),
    .A2(_00944_),
    .A3(_00946_),
    .A4(_00948_),
    .ZN(_00950_));
 BUF_X8 wire106 (.A(_01123_),
    .Z(net106));
 NAND2_X4 _05187_ (.A1(_00911_),
    .A2(net8),
    .ZN(_00952_));
 INV_X8 _05188_ (.A(net7),
    .ZN(_00953_));
 NAND3_X4 _05189_ (.A1(_00953_),
    .A2(net10),
    .A3(_00946_),
    .ZN(_00954_));
 BUF_X8 max_cap105 (.A(_01144_),
    .Z(net105));
 NOR2_X4 _05191_ (.A1(_00952_),
    .A2(_00954_),
    .ZN(_00956_));
 BUF_X8 max_cap104 (.A(net105),
    .Z(net104));
 BUF_X4 max_cap103 (.A(net105),
    .Z(net103));
 AOI221_X1 _05194_ (.A(_00943_),
    .B1(net266),
    .B2(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[12][0] ),
    .C1(net91),
    .C2(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[10][0] ),
    .ZN(_00959_));
 NAND2_X4 _05195_ (.A1(net1),
    .A2(net8),
    .ZN(_00960_));
 BUF_X4 wire102 (.A(net104),
    .Z(net102));
 OR3_X4 _05197_ (.A1(net7),
    .A2(net10),
    .A3(net9),
    .ZN(_00962_));
 BUF_X4 max_cap101 (.A(net104),
    .Z(net101));
 NOR2_X4 _05199_ (.A1(_00960_),
    .A2(_00962_),
    .ZN(_00964_));
 BUF_X4 max_cap100 (.A(net104),
    .Z(net100));
 BUF_X4 wire99 (.A(net105),
    .Z(net99));
 BUF_X8 max_cap98 (.A(net99),
    .Z(net98));
 BUF_X4 wire97 (.A(_01144_),
    .Z(net97));
 BUF_X16 max_cap96 (.A(_01149_),
    .Z(net96));
 NAND3_X4 _05205_ (.A1(_00953_),
    .A2(net10),
    .A3(net9),
    .ZN(_00970_));
 NOR2_X4 _05206_ (.A1(_00952_),
    .A2(_00970_),
    .ZN(_00971_));
 BUF_X16 max_cap95 (.A(net96),
    .Z(net95));
 BUF_X16 max_cap94 (.A(net95),
    .Z(net94));
 AOI22_X1 _05209_ (.A1(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[18][0] ),
    .A2(net264),
    .B1(net85),
    .B2(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[14][0] ),
    .ZN(_00974_));
 NOR4_X4 _05210_ (.A1(_00953_),
    .A2(net10),
    .A3(net9),
    .A4(_00948_),
    .ZN(_00975_));
 BUF_X16 max_cap93 (.A(net95),
    .Z(net93));
 BUF_X4 wire92 (.A(_01372_),
    .Z(net92));
 INV_X8 _05213_ (.A(net8),
    .ZN(_00978_));
 NAND2_X4 _05214_ (.A1(net1),
    .A2(_00978_),
    .ZN(_00979_));
 NAND3_X4 _05215_ (.A1(net7),
    .A2(_00944_),
    .A3(net9),
    .ZN(_00980_));
 NOR2_X4 _05216_ (.A1(_00979_),
    .A2(_00980_),
    .ZN(_00981_));
 BUF_X16 max_cap91 (.A(_00956_),
    .Z(net91));
 BUF_X16 max_length90 (.A(net91),
    .Z(net90));
 AOI22_X1 _05219_ (.A1(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[1][0] ),
    .A2(net258),
    .B1(net82),
    .B2(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[21][0] ),
    .ZN(_00984_));
 OR2_X4 _05220_ (.A1(net7),
    .A2(net10),
    .ZN(_00985_));
 NOR4_X4 _05221_ (.A1(_00911_),
    .A2(net8),
    .A3(_00946_),
    .A4(_00985_),
    .ZN(_00986_));
 BUF_X16 wire89 (.A(_00956_),
    .Z(net89));
 BUF_X16 max_cap88 (.A(_00971_),
    .Z(net88));
 NOR3_X4 _05224_ (.A1(net1),
    .A2(_00978_),
    .A3(_00962_),
    .ZN(_00989_));
 BUF_X16 max_cap87 (.A(_00971_),
    .Z(net87));
 AOI22_X1 _05226_ (.A1(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[20][0] ),
    .A2(net248),
    .B1(net243),
    .B2(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[2][0] ),
    .ZN(_00991_));
 NAND2_X4 _05227_ (.A1(net7),
    .A2(net10),
    .ZN(_00992_));
 NOR4_X4 _05228_ (.A1(net1),
    .A2(_00978_),
    .A3(net9),
    .A4(_00992_),
    .ZN(_00993_));
 BUF_X16 max_cap86 (.A(net87),
    .Z(net86));
 BUF_X16 max_cap85 (.A(net86),
    .Z(net85));
 NOR3_X4 _05231_ (.A1(_00946_),
    .A2(_00960_),
    .A3(_00985_),
    .ZN(_00996_));
 BUF_X16 max_cap84 (.A(_00981_),
    .Z(net84));
 AOI22_X1 _05233_ (.A1(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[11][0] ),
    .A2(net232),
    .B1(net223),
    .B2(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[22][0] ),
    .ZN(_00998_));
 NOR3_X4 _05234_ (.A1(net9),
    .A2(_00992_),
    .A3(_00948_),
    .ZN(_00999_));
 BUF_X16 max_cap83 (.A(net84),
    .Z(net83));
 BUF_X16 wire82 (.A(net84),
    .Z(net82));
 NOR4_X4 _05237_ (.A1(net7),
    .A2(_00944_),
    .A3(_00946_),
    .A4(_00960_),
    .ZN(_01002_));
 BUF_X16 max_cap81 (.A(_01019_),
    .Z(net81));
 AOI22_X1 _05239_ (.A1(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[9][0] ),
    .A2(net220),
    .B1(net207),
    .B2(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[30][0] ),
    .ZN(_01004_));
 NAND3_X4 _05240_ (.A1(net7),
    .A2(net10),
    .A3(net9),
    .ZN(_01005_));
 BUF_X16 max_length80 (.A(_01019_),
    .Z(net80));
 NOR2_X4 _05242_ (.A1(_01005_),
    .A2(_00948_),
    .ZN(_01007_));
 BUF_X16 max_length79 (.A(_01019_),
    .Z(net79));
 NOR4_X4 _05244_ (.A1(_00953_),
    .A2(net10),
    .A3(net9),
    .A4(_00960_),
    .ZN(_01009_));
 BUF_X16 max_cap78 (.A(net80),
    .Z(net78));
 AOI22_X1 _05246_ (.A1(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[13][0] ),
    .A2(net206),
    .B1(net197),
    .B2(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[19][0] ),
    .ZN(_01011_));
 AND4_X1 _05247_ (.A1(_00991_),
    .A2(_00998_),
    .A3(_01004_),
    .A4(_01011_),
    .ZN(_01012_));
 NAND4_X1 _05248_ (.A1(_00959_),
    .A2(_00974_),
    .A3(_00984_),
    .A4(_01012_),
    .ZN(_01013_));
 INV_X1 _05249_ (.A(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[3][0] ),
    .ZN(_01014_));
 NAND3_X4 _05250_ (.A1(net7),
    .A2(_00944_),
    .A3(_00946_),
    .ZN(_01015_));
 BUF_X16 max_cap77 (.A(_01032_),
    .Z(net77));
 INV_X1 _05252_ (.A(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[23][0] ),
    .ZN(_01017_));
 OAI33_X1 _05253_ (.A1(_01014_),
    .A2(_01015_),
    .A3(_00952_),
    .B1(_00980_),
    .B2(_00960_),
    .B3(_01017_),
    .ZN(_01018_));
 NOR2_X4 _05254_ (.A1(_01015_),
    .A2(_00979_),
    .ZN(_01019_));
 BUF_X16 max_cap76 (.A(_01032_),
    .Z(net76));
 NOR3_X4 _05256_ (.A1(net9),
    .A2(_00960_),
    .A3(_00992_),
    .ZN(_01021_));
 BUF_X16 max_cap75 (.A(net77),
    .Z(net75));
 AOI221_X1 _05258_ (.A(_01018_),
    .B1(net78),
    .B2(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[17][0] ),
    .C1(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[27][0] ),
    .C2(net191),
    .ZN(_01023_));
 INV_X1 _05259_ (.A(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[16][0] ),
    .ZN(_01024_));
 BUF_X16 max_cap74 (.A(_01059_),
    .Z(net74));
 NOR3_X4 _05261_ (.A1(net7),
    .A2(net10),
    .A3(net9),
    .ZN(_01026_));
 NAND3_X4 _05262_ (.A1(net1),
    .A2(_00978_),
    .A3(_01026_),
    .ZN(_01027_));
 BUF_X16 max_cap73 (.A(_01059_),
    .Z(net73));
 NAND3_X4 _05264_ (.A1(_00911_),
    .A2(net8),
    .A3(_00933_),
    .ZN(_01029_));
 INV_X1 _05265_ (.A(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[15][0] ),
    .ZN(_01030_));
 OAI22_X1 _05266_ (.A1(_01024_),
    .A2(_01027_),
    .B1(_01029_),
    .B2(_01030_),
    .ZN(_01031_));
 NOR2_X4 _05267_ (.A1(_00979_),
    .A2(_00970_),
    .ZN(_01032_));
 BUF_X16 max_cap72 (.A(net74),
    .Z(net72));
 NOR4_X4 _05269_ (.A1(net7),
    .A2(_00944_),
    .A3(net9),
    .A4(_00948_),
    .ZN(_01034_));
 BUF_X16 max_cap71 (.A(net74),
    .Z(net71));
 BUF_X16 max_cap70 (.A(_01076_),
    .Z(net70));
 AOI221_X1 _05272_ (.A(_01031_),
    .B1(net75),
    .B2(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[28][0] ),
    .C1(net183),
    .C2(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[8][0] ),
    .ZN(_01037_));
 NOR4_X4 _05273_ (.A1(net7),
    .A2(_00944_),
    .A3(net9),
    .A4(_00960_),
    .ZN(_01038_));
 BUF_X16 max_cap69 (.A(net70),
    .Z(net69));
 BUF_X16 max_cap68 (.A(_01076_),
    .Z(net68));
 BUF_X16 max_length67 (.A(net68),
    .Z(net67));
 NOR4_X4 _05277_ (.A1(net1),
    .A2(_00978_),
    .A3(_00946_),
    .A4(_00985_),
    .ZN(_01042_));
 BUF_X16 max_cap66 (.A(_01102_),
    .Z(net66));
 BUF_X16 max_cap65 (.A(net66),
    .Z(net65));
 AOI22_X1 _05280_ (.A1(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[26][0] ),
    .A2(net168),
    .B1(net164),
    .B2(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[6][0] ),
    .ZN(_01045_));
 NOR4_X4 _05281_ (.A1(_00911_),
    .A2(net8),
    .A3(net9),
    .A4(_00992_),
    .ZN(_01046_));
 BUF_X16 max_length64 (.A(net65),
    .Z(net64));
 BUF_X16 max_cap63 (.A(_01102_),
    .Z(net63));
 BUF_X4 output62 (.A(net62),
    .Z(valid_o));
 NOR3_X4 _05285_ (.A1(_00911_),
    .A2(net8),
    .A3(_01005_),
    .ZN(_01050_));
 BUF_X4 output61 (.A(net61),
    .Z(result_o[9]));
 BUF_X4 output60 (.A(net60),
    .Z(result_o[8]));
 AOI22_X1 _05288_ (.A1(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[25][0] ),
    .A2(net155),
    .B1(net145),
    .B2(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[29][0] ),
    .ZN(_01053_));
 AND2_X1 _05289_ (.A1(_01045_),
    .A2(_01053_),
    .ZN(_01054_));
 INV_X1 _05290_ (.A(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[7][0] ),
    .ZN(_01055_));
 OAI33_X1 _05291_ (.A1(_01055_),
    .A2(_00952_),
    .A3(_00980_),
    .B1(_00985_),
    .B2(_00948_),
    .B3(net9),
    .ZN(_01056_));
 NOR4_X4 _05292_ (.A1(_00953_),
    .A2(net10),
    .A3(_00946_),
    .A4(_00948_),
    .ZN(_01057_));
 BUF_X4 output59 (.A(net59),
    .Z(result_o[7]));
 NOR2_X4 _05294_ (.A1(_00979_),
    .A2(_00954_),
    .ZN(_01059_));
 BUF_X4 output58 (.A(net58),
    .Z(result_o[6]));
 BUF_X4 output57 (.A(net57),
    .Z(result_o[5]));
 AOI221_X1 _05297_ (.A(_01056_),
    .B1(net136),
    .B2(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[5][0] ),
    .C1(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[24][0] ),
    .C2(net72),
    .ZN(_01062_));
 NAND4_X1 _05298_ (.A1(_01023_),
    .A2(_01037_),
    .A3(_01054_),
    .A4(_01062_),
    .ZN(_01063_));
 NAND2_X4 _05299_ (.A1(_01026_),
    .A2(_00939_),
    .ZN(_01064_));
 BUF_X4 output56 (.A(net56),
    .Z(result_o[4]));
 BUF_X4 output55 (.A(net55),
    .Z(result_o[3]));
 BUF_X4 output54 (.A(net54),
    .Z(result_o[31]));
 OAI221_X1 _05303_ (.A(_00923_),
    .B1(_01013_),
    .B2(_01063_),
    .C1(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[0][0] ),
    .C2(_01064_),
    .ZN(_01068_));
 BUF_X4 output53 (.A(net53),
    .Z(result_o[30]));
 BUF_X4 output52 (.A(net52),
    .Z(result_o[2]));
 BUF_X4 output51 (.A(net51),
    .Z(result_o[29]));
 BUF_X4 output50 (.A(net50),
    .Z(result_o[28]));
 BUF_X4 output49 (.A(net49),
    .Z(result_o[27]));
 BUF_X4 output48 (.A(net48),
    .Z(result_o[26]));
 AOI22_X1 _05310_ (.A1(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[22][0] ),
    .A2(net223),
    .B1(net220),
    .B2(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[9][0] ),
    .ZN(_01075_));
 NOR2_X4 _05311_ (.A1(_00952_),
    .A2(_00980_),
    .ZN(_01076_));
 BUF_X4 output47 (.A(net47),
    .Z(result_o[25]));
 BUF_X4 output46 (.A(net46),
    .Z(result_o[24]));
 BUF_X4 output45 (.A(net45),
    .Z(result_o[23]));
 BUF_X4 output44 (.A(net44),
    .Z(result_o[22]));
 NOR3_X4 _05316_ (.A1(_00946_),
    .A2(_00985_),
    .A3(_00948_),
    .ZN(_01081_));
 BUF_X4 output43 (.A(net43),
    .Z(result_o[21]));
 BUF_X4 output42 (.A(net42),
    .Z(result_o[20]));
 AOI22_X1 _05319_ (.A1(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[7][0] ),
    .A2(net67),
    .B1(net125),
    .B2(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[4][0] ),
    .ZN(_01084_));
 BUF_X4 output41 (.A(net41),
    .Z(result_o[1]));
 BUF_X4 output40 (.A(net40),
    .Z(result_o[19]));
 BUF_X4 output39 (.A(net39),
    .Z(result_o[18]));
 BUF_X4 output38 (.A(net38),
    .Z(result_o[17]));
 BUF_X4 output37 (.A(net37),
    .Z(result_o[16]));
 BUF_X4 output36 (.A(net36),
    .Z(result_o[15]));
 AOI22_X1 _05326_ (.A1(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[12][0] ),
    .A2(net266),
    .B1(net258),
    .B2(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[1][0] ),
    .ZN(_01091_));
 BUF_X4 output35 (.A(net35),
    .Z(result_o[14]));
 BUF_X4 output34 (.A(net34),
    .Z(result_o[13]));
 BUF_X4 output33 (.A(net33),
    .Z(result_o[12]));
 AOI22_X1 _05330_ (.A1(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[17][0] ),
    .A2(net78),
    .B1(net191),
    .B2(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[27][0] ),
    .ZN(_01095_));
 NAND4_X1 _05331_ (.A1(_01075_),
    .A2(_01084_),
    .A3(_01091_),
    .A4(_01095_),
    .ZN(_01096_));
 NOR3_X4 _05332_ (.A1(_00911_),
    .A2(net8),
    .A3(_00962_),
    .ZN(_01097_));
 BUF_X4 output32 (.A(net32),
    .Z(result_o[11]));
 BUF_X4 output31 (.A(net31),
    .Z(result_o[10]));
 BUF_X4 output30 (.A(net30),
    .Z(result_o[0]));
 NAND2_X1 _05336_ (.A1(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[16][0] ),
    .A2(net119),
    .ZN(_01101_));
 NOR2_X4 _05337_ (.A1(_01015_),
    .A2(_00952_),
    .ZN(_01102_));
 BUF_X4 input29 (.A(we_i),
    .Z(net29));
 BUF_X1 input28 (.A(wdata_i[7]),
    .Z(net28));
 BUF_X1 input27 (.A(wdata_i[6]),
    .Z(net27));
 BUF_X1 input26 (.A(wdata_i[5]),
    .Z(net26));
 BUF_X1 input25 (.A(wdata_i[4]),
    .Z(net25));
 BUF_X1 input24 (.A(wdata_i[3]),
    .Z(net24));
 AOI22_X1 _05344_ (.A1(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[3][0] ),
    .A2(net65),
    .B1(net197),
    .B2(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[19][0] ),
    .ZN(_01109_));
 BUF_X1 input23 (.A(wdata_i[2]),
    .Z(net23));
 BUF_X1 input22 (.A(wdata_i[1]),
    .Z(net22));
 BUF_X1 input21 (.A(wdata_i[0]),
    .Z(net21));
 AOI22_X1 _05348_ (.A1(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[10][0] ),
    .A2(net91),
    .B1(net243),
    .B2(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[2][0] ),
    .ZN(_01113_));
 CLKBUF_X3 input20 (.A(waddr_i[8]),
    .Z(net20));
 BUF_X2 input19 (.A(waddr_i[7]),
    .Z(net19));
 BUF_X4 input18 (.A(waddr_i[6]),
    .Z(net18));
 AOI22_X1 _05352_ (.A1(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[25][0] ),
    .A2(net149),
    .B1(net248),
    .B2(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[20][0] ),
    .ZN(_01117_));
 NAND4_X1 _05353_ (.A1(_01101_),
    .A2(_01109_),
    .A3(_01113_),
    .A4(_01117_),
    .ZN(_01118_));
 NOR2_X4 _05354_ (.A1(_00962_),
    .A2(_00948_),
    .ZN(_01119_));
 BUF_X8 input17 (.A(waddr_i[5]),
    .Z(net17));
 NOR2_X4 _05356_ (.A1(_00911_),
    .A2(net8),
    .ZN(_01121_));
 AND2_X1 _05357_ (.A1(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[29][0] ),
    .A2(_01121_),
    .ZN(_01122_));
 NOR3_X4 _05358_ (.A1(net1),
    .A2(_00978_),
    .A3(_01005_),
    .ZN(_01123_));
 BUF_X4 input16 (.A(waddr_i[4]),
    .Z(net16));
 AOI221_X1 _05360_ (.A(net113),
    .B1(_01122_),
    .B2(_00933_),
    .C1(net109),
    .C2(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[15][0] ),
    .ZN(_01125_));
 BUF_X4 input15 (.A(waddr_i[3]),
    .Z(net15));
 BUF_X4 input14 (.A(waddr_i[2]),
    .Z(net14));
 BUF_X4 input13 (.A(waddr_i[1]),
    .Z(net13));
 BUF_X4 input12 (.A(waddr_i[0]),
    .Z(net12));
 BUF_X16 input11 (.A(rst_ni),
    .Z(net11));
 AOI22_X1 _05366_ (.A1(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[30][0] ),
    .A2(net207),
    .B1(net206),
    .B2(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[13][0] ),
    .ZN(_01131_));
 BUF_X16 input10 (.A(k_addr_i[3]),
    .Z(net10));
 BUF_X32 input9 (.A(k_addr_i[2]),
    .Z(net9));
 AOI22_X1 _05369_ (.A1(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[8][0] ),
    .A2(net183),
    .B1(net84),
    .B2(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[21][0] ),
    .ZN(_01134_));
 BUF_X16 input8 (.A(k_addr_i[1]),
    .Z(net8));
 BUF_X16 input7 (.A(k_addr_i[0]),
    .Z(net7));
 BUF_X4 input6 (.A(decoder_i),
    .Z(net6));
 BUF_X4 input5 (.A(c_addr_i[4]),
    .Z(net5));
 AOI22_X1 _05374_ (.A1(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[26][0] ),
    .A2(net168),
    .B1(net136),
    .B2(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[5][0] ),
    .ZN(_01139_));
 NAND4_X1 _05375_ (.A1(_01125_),
    .A2(_01131_),
    .A3(_01134_),
    .A4(_01139_),
    .ZN(_01140_));
 BUF_X8 input4 (.A(c_addr_i[3]),
    .Z(net4));
 BUF_X4 input3 (.A(c_addr_i[2]),
    .Z(net3));
 AOI22_X1 _05378_ (.A1(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[6][0] ),
    .A2(net160),
    .B1(net232),
    .B2(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[11][0] ),
    .ZN(_01143_));
 NOR4_X4 _05379_ (.A1(_00953_),
    .A2(net10),
    .A3(_00946_),
    .A4(_00960_),
    .ZN(_01144_));
 BUF_X4 input2 (.A(c_addr_i[1]),
    .Z(net2));
 BUF_X16 input1 (.A(c_addr_i[0]),
    .Z(net1));
 TAPCELL_X1 TAP_387 ();
 AOI22_X1 _05383_ (.A1(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[23][0] ),
    .A2(net98),
    .B1(net72),
    .B2(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[24][0] ),
    .ZN(_01148_));
 NOR2_X4 _05384_ (.A1(_00960_),
    .A2(_01005_),
    .ZN(_01149_));
 TAPCELL_X1 TAP_386 ();
 TAPCELL_X1 TAP_385 ();
 TAPCELL_X1 TAP_384 ();
 TAPCELL_X1 TAP_383 ();
 TAPCELL_X1 TAP_382 ();
 AOI22_X1 _05390_ (.A1(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[31][0] ),
    .A2(_01149_),
    .B1(net264),
    .B2(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[18][0] ),
    .ZN(_01155_));
 TAPCELL_X1 TAP_381 ();
 TAPCELL_X1 TAP_380 ();
 TAPCELL_X1 TAP_379 ();
 TAPCELL_X1 TAP_378 ();
 AOI22_X1 _05395_ (.A1(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[28][0] ),
    .A2(net75),
    .B1(net86),
    .B2(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[14][0] ),
    .ZN(_01160_));
 NAND4_X1 _05396_ (.A1(_01143_),
    .A2(_01148_),
    .A3(_01155_),
    .A4(_01160_),
    .ZN(_01161_));
 NOR4_X2 _05397_ (.A1(_01096_),
    .A2(_01118_),
    .A3(_01140_),
    .A4(_01161_),
    .ZN(_01162_));
 NAND2_X4 _05398_ (.A1(net4),
    .A2(net5),
    .ZN(_01163_));
 NOR3_X4 _05399_ (.A1(net2),
    .A2(net3),
    .A3(_01163_),
    .ZN(_01164_));
 TAPCELL_X1 TAP_377 ();
 OAI21_X1 _05401_ (.A(_01164_),
    .B1(_01064_),
    .B2(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[0][0] ),
    .ZN(_01166_));
 OAI21_X1 _05402_ (.A(_01068_),
    .B1(_01162_),
    .B2(_01166_),
    .ZN(_01167_));
 NAND2_X4 _05403_ (.A1(net4),
    .A2(_00920_),
    .ZN(_01168_));
 NOR3_X4 _05404_ (.A1(net2),
    .A2(net3),
    .A3(_01168_),
    .ZN(_01169_));
 INV_X1 _05405_ (.A(_01169_),
    .ZN(_01170_));
 TAPCELL_X1 TAP_376 ();
 TAPCELL_X1 TAP_375 ();
 TAPCELL_X1 TAP_374 ();
 AOI22_X1 _05409_ (.A1(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[27][0] ),
    .A2(net190),
    .B1(net113),
    .B2(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[0][0] ),
    .ZN(_01174_));
 TAPCELL_X1 TAP_373 ();
 TAPCELL_X1 TAP_372 ();
 AOI22_X1 _05412_ (.A1(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[24][0] ),
    .A2(net74),
    .B1(net249),
    .B2(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[20][0] ),
    .ZN(_01177_));
 AOI22_X1 _05413_ (.A1(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[25][0] ),
    .A2(net155),
    .B1(net195),
    .B2(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[19][0] ),
    .ZN(_01178_));
 TAPCELL_X1 TAP_371 ();
 AOI22_X1 _05415_ (.A1(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[3][0] ),
    .A2(net64),
    .B1(net137),
    .B2(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[5][0] ),
    .ZN(_01180_));
 NAND4_X1 _05416_ (.A1(_01174_),
    .A2(_01177_),
    .A3(_01178_),
    .A4(_01180_),
    .ZN(_01181_));
 TAPCELL_X1 TAP_370 ();
 AOI22_X1 _05418_ (.A1(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[17][0] ),
    .A2(net80),
    .B1(net75),
    .B2(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[28][0] ),
    .ZN(_01183_));
 AOI22_X1 _05419_ (.A1(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[23][0] ),
    .A2(net103),
    .B1(net82),
    .B2(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[21][0] ),
    .ZN(_01184_));
 TAPCELL_X1 TAP_369 ();
 TAPCELL_X1 TAP_368 ();
 TAPCELL_X1 TAP_367 ();
 TAPCELL_X1 TAP_366 ();
 TAPCELL_X1 TAP_365 ();
 AOI22_X1 _05425_ (.A1(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[16][0] ),
    .A2(net118),
    .B1(net161),
    .B2(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[6][0] ),
    .ZN(_01190_));
 TAPCELL_X1 TAP_364 ();
 TAPCELL_X1 TAP_363 ();
 TAPCELL_X1 TAP_362 ();
 AOI22_X2 _05429_ (.A1(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[31][0] ),
    .A2(net96),
    .B1(net205),
    .B2(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[13][0] ),
    .ZN(_01194_));
 NAND4_X2 _05430_ (.A1(_01183_),
    .A2(_01184_),
    .A3(_01190_),
    .A4(_01194_),
    .ZN(_01195_));
 TAPCELL_X1 TAP_361 ();
 AOI22_X1 _05432_ (.A1(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[11][0] ),
    .A2(net235),
    .B1(net219),
    .B2(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[9][0] ),
    .ZN(_01197_));
 TAPCELL_X1 TAP_360 ();
 AOI22_X1 _05434_ (.A1(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[8][0] ),
    .A2(net184),
    .B1(net124),
    .B2(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[4][0] ),
    .ZN(_01199_));
 AND2_X1 _05435_ (.A1(_01197_),
    .A2(_01199_),
    .ZN(_01200_));
 INV_X1 _05436_ (.A(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[26][0] ),
    .ZN(_01201_));
 TAPCELL_X1 TAP_359 ();
 NAND4_X4 _05438_ (.A1(_00953_),
    .A2(net10),
    .A3(_00946_),
    .A4(_00926_),
    .ZN(_01203_));
 NAND4_X4 _05439_ (.A1(_00953_),
    .A2(net10),
    .A3(net9),
    .A4(_00926_),
    .ZN(_01204_));
 INV_X1 _05440_ (.A(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[30][0] ),
    .ZN(_01205_));
 OAI22_X1 _05441_ (.A1(_01201_),
    .A2(_01203_),
    .B1(_01204_),
    .B2(_01205_),
    .ZN(_01206_));
 TAPCELL_X1 TAP_358 ();
 AOI221_X1 _05443_ (.A(_01206_),
    .B1(net85),
    .B2(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[14][0] ),
    .C1(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[18][0] ),
    .C2(net265),
    .ZN(_01208_));
 INV_X1 _05444_ (.A(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[1][0] ),
    .ZN(_01209_));
 NAND4_X4 _05445_ (.A1(net7),
    .A2(_00944_),
    .A3(_00946_),
    .A4(_00939_),
    .ZN(_01210_));
 NAND3_X4 _05446_ (.A1(_00911_),
    .A2(net8),
    .A3(_01026_),
    .ZN(_01211_));
 INV_X1 _05447_ (.A(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[2][0] ),
    .ZN(_01212_));
 OAI22_X1 _05448_ (.A1(_01209_),
    .A2(_01210_),
    .B1(_01211_),
    .B2(_01212_),
    .ZN(_01213_));
 AOI221_X1 _05449_ (.A(_01213_),
    .B1(net67),
    .B2(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[7][0] ),
    .C1(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[12][0] ),
    .C2(net271),
    .ZN(_01214_));
 INV_X1 _05450_ (.A(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[15][0] ),
    .ZN(_01215_));
 NAND3_X4 _05451_ (.A1(net9),
    .A2(_00926_),
    .A3(_00937_),
    .ZN(_01216_));
 INV_X1 _05452_ (.A(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[22][0] ),
    .ZN(_01217_));
 OAI22_X1 _05453_ (.A1(_01215_),
    .A2(_01029_),
    .B1(_01216_),
    .B2(_01217_),
    .ZN(_01218_));
 TAPCELL_X1 TAP_357 ();
 AOI221_X1 _05455_ (.A(_01218_),
    .B1(net90),
    .B2(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[10][0] ),
    .C1(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[29][0] ),
    .C2(net145),
    .ZN(_01220_));
 NAND4_X1 _05456_ (.A1(_01200_),
    .A2(_01208_),
    .A3(_01214_),
    .A4(_01220_),
    .ZN(_01221_));
 NOR3_X1 _05457_ (.A1(_01181_),
    .A2(_01195_),
    .A3(_01221_),
    .ZN(_01222_));
 TAPCELL_X1 TAP_356 ();
 TAPCELL_X1 TAP_355 ();
 AOI22_X1 _05460_ (.A1(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[28][0] ),
    .A2(net76),
    .B1(net144),
    .B2(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[29][0] ),
    .ZN(_01225_));
 TAPCELL_X1 TAP_354 ();
 TAPCELL_X1 TAP_353 ();
 TAPCELL_X1 TAP_352 ();
 TAPCELL_X1 TAP_351 ();
 TAPCELL_X1 TAP_350 ();
 AOI22_X1 _05466_ (.A1(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[7][0] ),
    .A2(net69),
    .B1(net126),
    .B2(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[4][0] ),
    .ZN(_01231_));
 TAPCELL_X1 TAP_349 ();
 TAPCELL_X1 TAP_348 ();
 TAPCELL_X1 TAP_347 ();
 TAPCELL_X1 TAP_346 ();
 AOI22_X1 _05471_ (.A1(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[23][0] ),
    .A2(net102),
    .B1(net196),
    .B2(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[19][0] ),
    .ZN(_01236_));
 TAPCELL_X1 TAP_345 ();
 TAPCELL_X1 TAP_344 ();
 TAPCELL_X1 TAP_343 ();
 AOI22_X2 _05475_ (.A1(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[15][0] ),
    .A2(net108),
    .B1(net245),
    .B2(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[20][0] ),
    .ZN(_01240_));
 NAND4_X2 _05476_ (.A1(_01225_),
    .A2(_01231_),
    .A3(_01236_),
    .A4(_01240_),
    .ZN(_01241_));
 TAPCELL_X1 TAP_342 ();
 TAPCELL_X1 TAP_341 ();
 TAPCELL_X1 TAP_340 ();
 TAPCELL_X1 TAP_339 ();
 AOI22_X1 _05481_ (.A1(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[26][0] ),
    .A2(net174),
    .B1(net263),
    .B2(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[18][0] ),
    .ZN(_01246_));
 TAPCELL_X1 TAP_338 ();
 TAPCELL_X1 TAP_337 ();
 TAPCELL_X1 TAP_336 ();
 AOI22_X1 _05485_ (.A1(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[10][0] ),
    .A2(_00956_),
    .B1(net87),
    .B2(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[14][0] ),
    .ZN(_01250_));
 TAPCELL_X1 TAP_335 ();
 TAPCELL_X1 TAP_334 ();
 TAPCELL_X1 TAP_333 ();
 TAPCELL_X1 TAP_332 ();
 AOI22_X1 _05490_ (.A1(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[24][0] ),
    .A2(net71),
    .B1(net213),
    .B2(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[30][0] ),
    .ZN(_01255_));
 TAPCELL_X1 TAP_331 ();
 TAPCELL_X1 TAP_330 ();
 TAPCELL_X1 TAP_329 ();
 AOI21_X1 _05494_ (.A(net114),
    .B1(net217),
    .B2(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[9][0] ),
    .ZN(_01259_));
 NAND4_X2 _05495_ (.A1(_01246_),
    .A2(_01250_),
    .A3(_01255_),
    .A4(_01259_),
    .ZN(_01260_));
 TAPCELL_X1 TAP_328 ();
 TAPCELL_X1 TAP_327 ();
 AOI22_X1 _05498_ (.A1(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[16][0] ),
    .A2(net120),
    .B1(net83),
    .B2(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[21][0] ),
    .ZN(_01263_));
 TAPCELL_X1 TAP_326 ();
 TAPCELL_X1 TAP_325 ();
 TAPCELL_X1 TAP_324 ();
 TAPCELL_X1 TAP_323 ();
 AOI22_X1 _05503_ (.A1(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[3][0] ),
    .A2(net66),
    .B1(net229),
    .B2(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[11][0] ),
    .ZN(_01268_));
 TAPCELL_X1 TAP_322 ();
 TAPCELL_X1 TAP_321 ();
 TAPCELL_X1 TAP_320 ();
 TAPCELL_X1 TAP_319 ();
 AOI22_X1 _05508_ (.A1(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[27][0] ),
    .A2(net188),
    .B1(net238),
    .B2(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[2][0] ),
    .ZN(_01273_));
 TAPCELL_X1 TAP_318 ();
 AOI22_X2 _05510_ (.A1(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[22][0] ),
    .A2(net222),
    .B1(net203),
    .B2(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[13][0] ),
    .ZN(_01275_));
 NAND4_X2 _05511_ (.A1(_01263_),
    .A2(_01268_),
    .A3(_01273_),
    .A4(_01275_),
    .ZN(_01276_));
 TAPCELL_X1 TAP_317 ();
 TAPCELL_X1 TAP_316 ();
 TAPCELL_X1 TAP_315 ();
 AOI22_X1 _05515_ (.A1(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[6][0] ),
    .A2(net158),
    .B1(net134),
    .B2(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[5][0] ),
    .ZN(_01280_));
 TAPCELL_X1 TAP_314 ();
 TAPCELL_X1 TAP_313 ();
 TAPCELL_X1 TAP_312 ();
 AOI22_X1 _05519_ (.A1(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[25][0] ),
    .A2(net152),
    .B1(net93),
    .B2(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[31][0] ),
    .ZN(_01284_));
 TAPCELL_X1 TAP_311 ();
 TAPCELL_X1 TAP_310 ();
 TAPCELL_X1 PHY_309 ();
 AOI22_X2 _05523_ (.A1(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[17][0] ),
    .A2(net79),
    .B1(net254),
    .B2(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[1][0] ),
    .ZN(_01288_));
 TAPCELL_X1 PHY_308 ();
 TAPCELL_X1 PHY_307 ();
 TAPCELL_X1 PHY_306 ();
 AOI22_X2 _05527_ (.A1(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[8][0] ),
    .A2(net178),
    .B1(net268),
    .B2(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[12][0] ),
    .ZN(_01292_));
 NAND4_X2 _05528_ (.A1(_01280_),
    .A2(_01284_),
    .A3(_01288_),
    .A4(_01292_),
    .ZN(_01293_));
 NOR4_X4 _05529_ (.A1(_01241_),
    .A2(_01260_),
    .A3(_01276_),
    .A4(_01293_),
    .ZN(_01294_));
 NOR2_X4 _05530_ (.A1(_00921_),
    .A2(_01168_),
    .ZN(_01295_));
 TAPCELL_X1 PHY_305 ();
 TAPCELL_X1 PHY_304 ();
 OAI21_X1 _05533_ (.A(_01295_),
    .B1(net130),
    .B2(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[0][0] ),
    .ZN(_01298_));
 OAI22_X1 _05534_ (.A1(_01170_),
    .A2(_01222_),
    .B1(_01294_),
    .B2(_01298_),
    .ZN(_01299_));
 TAPCELL_X1 PHY_303 ();
 AOI22_X1 _05536_ (.A1(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[28][0] ),
    .A2(net75),
    .B1(net85),
    .B2(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[14][0] ),
    .ZN(_01301_));
 TAPCELL_X1 PHY_302 ();
 AOI22_X1 _05538_ (.A1(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[5][0] ),
    .A2(net138),
    .B1(net241),
    .B2(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[2][0] ),
    .ZN(_01303_));
 TAPCELL_X1 PHY_301 ();
 AOI22_X1 _05540_ (.A1(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[8][0] ),
    .A2(net184),
    .B1(net72),
    .B2(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[24][0] ),
    .ZN(_01305_));
 TAPCELL_X1 PHY_300 ();
 TAPCELL_X1 PHY_299 ();
 TAPCELL_X1 PHY_298 ();
 AOI22_X1 _05544_ (.A1(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[12][0] ),
    .A2(net270),
    .B1(net257),
    .B2(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[1][0] ),
    .ZN(_01309_));
 NAND4_X1 _05545_ (.A1(_01301_),
    .A2(_01303_),
    .A3(_01305_),
    .A4(_01309_),
    .ZN(_01310_));
 TAPCELL_X1 PHY_297 ();
 AOI22_X1 _05547_ (.A1(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[11][0] ),
    .A2(net235),
    .B1(net225),
    .B2(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[22][0] ),
    .ZN(_01312_));
 TAPCELL_X1 PHY_296 ();
 TAPCELL_X1 PHY_295 ();
 AOI22_X1 _05550_ (.A1(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[17][0] ),
    .A2(net80),
    .B1(net169),
    .B2(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[26][0] ),
    .ZN(_01315_));
 TAPCELL_X1 PHY_294 ();
 TAPCELL_X1 PHY_293 ();
 TAPCELL_X1 PHY_292 ();
 AOI22_X1 _05554_ (.A1(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[29][0] ),
    .A2(net143),
    .B1(net96),
    .B2(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[31][0] ),
    .ZN(_01319_));
 AOI21_X1 _05555_ (.A(net113),
    .B1(net197),
    .B2(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[19][0] ),
    .ZN(_01320_));
 NAND4_X1 _05556_ (.A1(_01312_),
    .A2(_01315_),
    .A3(_01319_),
    .A4(_01320_),
    .ZN(_01321_));
 TAPCELL_X1 PHY_291 ();
 AOI22_X1 _05558_ (.A1(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[10][0] ),
    .A2(net91),
    .B1(net210),
    .B2(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[30][0] ),
    .ZN(_01323_));
 TAPCELL_X1 PHY_290 ();
 TAPCELL_X1 PHY_289 ();
 AOI22_X1 _05561_ (.A1(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[3][0] ),
    .A2(net64),
    .B1(net118),
    .B2(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[16][0] ),
    .ZN(_01326_));
 TAPCELL_X1 PHY_288 ();
 TAPCELL_X1 PHY_287 ();
 TAPCELL_X1 PHY_286 ();
 AOI22_X1 _05565_ (.A1(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[15][0] ),
    .A2(net106),
    .B1(net219),
    .B2(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[9][0] ),
    .ZN(_01330_));
 TAPCELL_X1 PHY_285 ();
 TAPCELL_X1 PHY_284 ();
 AOI22_X1 _05568_ (.A1(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[6][0] ),
    .A2(net161),
    .B1(net82),
    .B2(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[21][0] ),
    .ZN(_01333_));
 NAND4_X2 _05569_ (.A1(_01323_),
    .A2(_01326_),
    .A3(_01330_),
    .A4(_01333_),
    .ZN(_01334_));
 TAPCELL_X1 PHY_283 ();
 TAPCELL_X1 PHY_282 ();
 TAPCELL_X1 PHY_281 ();
 TAPCELL_X1 PHY_280 ();
 AOI22_X1 _05574_ (.A1(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[23][0] ),
    .A2(net103),
    .B1(net125),
    .B2(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[4][0] ),
    .ZN(_01339_));
 TAPCELL_X1 PHY_279 ();
 TAPCELL_X1 PHY_278 ();
 AOI22_X1 _05577_ (.A1(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[27][0] ),
    .A2(net189),
    .B1(net247),
    .B2(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[20][0] ),
    .ZN(_01342_));
 TAPCELL_X1 PHY_277 ();
 AOI22_X1 _05579_ (.A1(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[7][0] ),
    .A2(net67),
    .B1(net264),
    .B2(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[18][0] ),
    .ZN(_01344_));
 TAPCELL_X1 PHY_276 ();
 AOI22_X2 _05581_ (.A1(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[25][0] ),
    .A2(net154),
    .B1(net205),
    .B2(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[13][0] ),
    .ZN(_01346_));
 NAND4_X2 _05582_ (.A1(_01339_),
    .A2(_01342_),
    .A3(_01344_),
    .A4(_01346_),
    .ZN(_01347_));
 NOR4_X2 _05583_ (.A1(_01310_),
    .A2(_01321_),
    .A3(_01334_),
    .A4(_01347_),
    .ZN(_01348_));
 NAND2_X4 _05584_ (.A1(net2),
    .A2(net3),
    .ZN(_01349_));
 NOR2_X4 _05585_ (.A1(_01168_),
    .A2(_01349_),
    .ZN(_01350_));
 OAI21_X1 _05586_ (.A(_01350_),
    .B1(net130),
    .B2(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[0][0] ),
    .ZN(_01351_));
 TAPCELL_X1 PHY_275 ();
 TAPCELL_X1 PHY_274 ();
 TAPCELL_X1 PHY_273 ();
 TAPCELL_X1 PHY_272 ();
 AOI22_X1 _05591_ (.A1(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[25][0] ),
    .A2(net152),
    .B1(net83),
    .B2(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[21][0] ),
    .ZN(_01356_));
 TAPCELL_X1 PHY_271 ();
 AOI22_X1 _05593_ (.A1(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[15][0] ),
    .A2(net107),
    .B1(net217),
    .B2(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[9][0] ),
    .ZN(_01358_));
 TAPCELL_X1 PHY_270 ();
 AOI22_X1 _05595_ (.A1(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[3][0] ),
    .A2(net66),
    .B1(net71),
    .B2(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[24][0] ),
    .ZN(_01360_));
 TAPCELL_X1 PHY_269 ();
 TAPCELL_X1 PHY_268 ();
 AOI22_X1 _05598_ (.A1(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[26][0] ),
    .A2(net173),
    .B1(net68),
    .B2(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[7][0] ),
    .ZN(_01363_));
 NAND4_X1 _05599_ (.A1(_01356_),
    .A2(_01358_),
    .A3(_01360_),
    .A4(_01363_),
    .ZN(_01364_));
 TAPCELL_X1 PHY_267 ();
 AOI22_X1 _05601_ (.A1(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[28][0] ),
    .A2(net76),
    .B1(net222),
    .B2(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[22][0] ),
    .ZN(_01366_));
 TAPCELL_X1 PHY_266 ();
 TAPCELL_X1 PHY_265 ();
 TAPCELL_X1 PHY_264 ();
 AOI22_X1 _05605_ (.A1(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[2][0] ),
    .A2(net240),
    .B1(net193),
    .B2(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[19][0] ),
    .ZN(_01370_));
 TAPCELL_X1 PHY_263 ();
 NOR4_X2 _05607_ (.A1(net1),
    .A2(net7),
    .A3(_00944_),
    .A4(_00946_),
    .ZN(_01372_));
 TAPCELL_X1 PHY_262 ();
 MUX2_X1 _05609_ (.A(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[12][0] ),
    .B(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[14][0] ),
    .S(net8),
    .Z(_01374_));
 TAPCELL_X1 PHY_261 ();
 AOI221_X1 _05611_ (.A(net114),
    .B1(net92),
    .B2(_01374_),
    .C1(net254),
    .C2(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[1][0] ),
    .ZN(_01376_));
 NAND3_X1 _05612_ (.A1(_01366_),
    .A2(_01370_),
    .A3(_01376_),
    .ZN(_01377_));
 TAPCELL_X1 PHY_260 ();
 TAPCELL_X1 PHY_259 ();
 AOI22_X1 _05615_ (.A1(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[8][0] ),
    .A2(net180),
    .B1(net123),
    .B2(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[4][0] ),
    .ZN(_01380_));
 TAPCELL_X1 PHY_258 ();
 AOI22_X1 _05617_ (.A1(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[17][0] ),
    .A2(net79),
    .B1(net90),
    .B2(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[10][0] ),
    .ZN(_01382_));
 TAPCELL_X1 PHY_257 ();
 TAPCELL_X1 PHY_256 ();
 AOI22_X1 _05620_ (.A1(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[6][0] ),
    .A2(net162),
    .B1(net144),
    .B2(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[29][0] ),
    .ZN(_01385_));
 TAPCELL_X1 PHY_255 ();
 AOI22_X2 _05622_ (.A1(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[18][0] ),
    .A2(net263),
    .B1(net204),
    .B2(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[13][0] ),
    .ZN(_01387_));
 NAND4_X2 _05623_ (.A1(_01380_),
    .A2(_01382_),
    .A3(_01385_),
    .A4(_01387_),
    .ZN(_01388_));
 TAPCELL_X1 PHY_254 ();
 TAPCELL_X1 PHY_253 ();
 AOI22_X1 _05626_ (.A1(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[20][0] ),
    .A2(net250),
    .B1(net208),
    .B2(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[30][0] ),
    .ZN(_01391_));
 TAPCELL_X1 PHY_252 ();
 TAPCELL_X1 PHY_251 ();
 AOI22_X1 _05629_ (.A1(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[27][0] ),
    .A2(net188),
    .B1(net116),
    .B2(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[16][0] ),
    .ZN(_01394_));
 TAPCELL_X1 PHY_250 ();
 AOI22_X1 _05631_ (.A1(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[23][0] ),
    .A2(net100),
    .B1(net93),
    .B2(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[31][0] ),
    .ZN(_01396_));
 TAPCELL_X1 PHY_249 ();
 AOI22_X2 _05633_ (.A1(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[5][0] ),
    .A2(net131),
    .B1(net233),
    .B2(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[11][0] ),
    .ZN(_01398_));
 NAND4_X2 _05634_ (.A1(_01391_),
    .A2(_01394_),
    .A3(_01396_),
    .A4(_01398_),
    .ZN(_01399_));
 NOR4_X2 _05635_ (.A1(_01364_),
    .A2(_01377_),
    .A3(_01388_),
    .A4(_01399_),
    .ZN(_01400_));
 NOR2_X2 _05636_ (.A1(_00922_),
    .A2(_01349_),
    .ZN(_01401_));
 TAPCELL_X1 PHY_248 ();
 TAPCELL_X1 PHY_247 ();
 OAI21_X1 _05639_ (.A(_01401_),
    .B1(net130),
    .B2(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[0][0] ),
    .ZN(_01404_));
 OAI22_X1 _05640_ (.A1(_01348_),
    .A2(_01351_),
    .B1(_01400_),
    .B2(_01404_),
    .ZN(_01405_));
 NAND4_X4 _05641_ (.A1(_00914_),
    .A2(_00916_),
    .A3(_00918_),
    .A4(_00920_),
    .ZN(_01406_));
 NAND2_X4 _05642_ (.A1(_00914_),
    .A2(net3),
    .ZN(_01407_));
 NOR2_X2 _05643_ (.A1(_01168_),
    .A2(_01407_),
    .ZN(_01408_));
 TAPCELL_X1 PHY_246 ();
 OAI21_X1 _05645_ (.A(_01408_),
    .B1(net130),
    .B2(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[0][0] ),
    .ZN(_01410_));
 INV_X1 _05646_ (.A(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[15][0] ),
    .ZN(_01411_));
 INV_X1 _05647_ (.A(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[2][0] ),
    .ZN(_01412_));
 OAI22_X1 _05648_ (.A1(_01411_),
    .A2(_01029_),
    .B1(_01211_),
    .B2(_01412_),
    .ZN(_01413_));
 TAPCELL_X1 PHY_245 ();
 AOI221_X1 _05650_ (.A(_01413_),
    .B1(_01076_),
    .B2(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[7][0] ),
    .C1(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[27][0] ),
    .C2(net192),
    .ZN(_01415_));
 INV_X1 _05651_ (.A(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[23][0] ),
    .ZN(_01416_));
 NAND4_X4 _05652_ (.A1(net7),
    .A2(_00944_),
    .A3(net9),
    .A4(_00926_),
    .ZN(_01417_));
 AND2_X4 _05653_ (.A1(net7),
    .A2(net10),
    .ZN(_01418_));
 TAPCELL_X1 PHY_244 ();
 NAND3_X4 _05655_ (.A1(_00946_),
    .A2(_01418_),
    .A3(_00939_),
    .ZN(_01420_));
 INV_X1 _05656_ (.A(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[9][0] ),
    .ZN(_01421_));
 OAI22_X1 _05657_ (.A1(_01416_),
    .A2(_01417_),
    .B1(_01420_),
    .B2(_01421_),
    .ZN(_01422_));
 AOI221_X1 _05658_ (.A(_01422_),
    .B1(_01034_),
    .B2(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[8][0] ),
    .C1(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[14][0] ),
    .C2(net87),
    .ZN(_01423_));
 INV_X1 _05659_ (.A(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[29][0] ),
    .ZN(_01424_));
 NAND3_X4 _05660_ (.A1(net1),
    .A2(_00978_),
    .A3(_00933_),
    .ZN(_01425_));
 NAND4_X4 _05661_ (.A1(_00953_),
    .A2(net10),
    .A3(net9),
    .A4(_00939_),
    .ZN(_01426_));
 INV_X1 _05662_ (.A(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[12][0] ),
    .ZN(_01427_));
 OAI22_X1 _05663_ (.A1(_01424_),
    .A2(_01425_),
    .B1(_01426_),
    .B2(_01427_),
    .ZN(_01428_));
 AOI221_X1 _05664_ (.A(_01428_),
    .B1(net128),
    .B2(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[4][0] ),
    .C1(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[24][0] ),
    .C2(net73),
    .ZN(_01429_));
 INV_X1 _05665_ (.A(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[28][0] ),
    .ZN(_01430_));
 TAPCELL_X1 PHY_243 ();
 OAI33_X1 _05667_ (.A1(_01430_),
    .A2(_00979_),
    .A3(_00970_),
    .B1(_00948_),
    .B2(_00985_),
    .B3(net9),
    .ZN(_01432_));
 AOI221_X1 _05668_ (.A(_01432_),
    .B1(net225),
    .B2(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[22][0] ),
    .C1(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[30][0] ),
    .C2(net211),
    .ZN(_01433_));
 NAND4_X1 _05669_ (.A1(_01415_),
    .A2(_01423_),
    .A3(_01429_),
    .A4(_01433_),
    .ZN(_01434_));
 AOI22_X1 _05670_ (.A1(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[6][0] ),
    .A2(net156),
    .B1(net206),
    .B2(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[13][0] ),
    .ZN(_01435_));
 TAPCELL_X1 PHY_242 ();
 AOI22_X1 _05672_ (.A1(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[26][0] ),
    .A2(net171),
    .B1(net253),
    .B2(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[1][0] ),
    .ZN(_01437_));
 TAPCELL_X1 PHY_241 ();
 TAPCELL_X1 PHY_240 ();
 AOI22_X1 _05675_ (.A1(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[25][0] ),
    .A2(net150),
    .B1(net139),
    .B2(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[5][0] ),
    .ZN(_01440_));
 TAPCELL_X1 PHY_239 ();
 TAPCELL_X1 PHY_238 ();
 AOI22_X2 _05678_ (.A1(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[10][0] ),
    .A2(net89),
    .B1(net201),
    .B2(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[19][0] ),
    .ZN(_01443_));
 NAND4_X2 _05679_ (.A1(_01435_),
    .A2(_01437_),
    .A3(_01440_),
    .A4(_01443_),
    .ZN(_01444_));
 TAPCELL_X1 PHY_237 ();
 AOI22_X1 _05681_ (.A1(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[18][0] ),
    .A2(net264),
    .B1(net248),
    .B2(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[20][0] ),
    .ZN(_01446_));
 TAPCELL_X1 PHY_236 ();
 AOI22_X1 _05683_ (.A1(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[17][0] ),
    .A2(net78),
    .B1(net84),
    .B2(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[21][0] ),
    .ZN(_01448_));
 TAPCELL_X1 PHY_235 ();
 TAPCELL_X1 PHY_234 ();
 TAPCELL_X1 PHY_233 ();
 AOI22_X1 _05687_ (.A1(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[3][0] ),
    .A2(net65),
    .B1(net237),
    .B2(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[11][0] ),
    .ZN(_01452_));
 TAPCELL_X1 PHY_232 ();
 AOI22_X1 _05689_ (.A1(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[16][0] ),
    .A2(net119),
    .B1(_01149_),
    .B2(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[31][0] ),
    .ZN(_01454_));
 NAND4_X1 _05690_ (.A1(_01446_),
    .A2(_01448_),
    .A3(_01452_),
    .A4(_01454_),
    .ZN(_01455_));
 NOR3_X1 _05691_ (.A1(_01434_),
    .A2(_01444_),
    .A3(_01455_),
    .ZN(_01456_));
 OAI21_X1 _05692_ (.A(_01406_),
    .B1(_01410_),
    .B2(_01456_),
    .ZN(_01457_));
 NOR4_X1 _05693_ (.A1(_01167_),
    .A2(_01299_),
    .A3(_01405_),
    .A4(_01457_),
    .ZN(_01458_));
 INV_X1 _05694_ (.A(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[23][0] ),
    .ZN(_01459_));
 INV_X1 _05695_ (.A(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[2][0] ),
    .ZN(_01460_));
 OAI22_X1 _05696_ (.A1(_01459_),
    .A2(_01417_),
    .B1(_01211_),
    .B2(_01460_),
    .ZN(_01461_));
 TAPCELL_X1 PHY_231 ();
 AOI221_X1 _05698_ (.A(_01461_),
    .B1(_00964_),
    .B2(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[18][0] ),
    .C1(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[21][0] ),
    .C2(_00981_),
    .ZN(_01463_));
 TAPCELL_X1 PHY_230 ();
 AOI22_X1 _05700_ (.A1(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[12][0] ),
    .A2(net274),
    .B1(net215),
    .B2(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[30][0] ),
    .ZN(_01465_));
 TAPCELL_X1 PHY_229 ();
 AOI22_X1 _05702_ (.A1(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[8][0] ),
    .A2(net176),
    .B1(net156),
    .B2(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[6][0] ),
    .ZN(_01467_));
 AND2_X1 _05703_ (.A1(_01465_),
    .A2(_01467_),
    .ZN(_01468_));
 INV_X1 _05704_ (.A(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[25][0] ),
    .ZN(_01469_));
 NAND4_X4 _05705_ (.A1(net1),
    .A2(_00978_),
    .A3(_00946_),
    .A4(_01418_),
    .ZN(_01470_));
 INV_X1 _05706_ (.A(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[9][0] ),
    .ZN(_01471_));
 OAI22_X1 _05707_ (.A1(_01469_),
    .A2(_01470_),
    .B1(_01420_),
    .B2(_01471_),
    .ZN(_01472_));
 TAPCELL_X1 PHY_228 ();
 AOI221_X1 _05709_ (.A(_01472_),
    .B1(net129),
    .B2(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[4][0] ),
    .C1(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[7][0] ),
    .C2(net70),
    .ZN(_01474_));
 INV_X1 _05710_ (.A(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[26][0] ),
    .ZN(_01475_));
 OAI21_X1 _05711_ (.A(_01064_),
    .B1(_01203_),
    .B2(_01475_),
    .ZN(_01476_));
 TAPCELL_X1 PHY_227 ();
 TAPCELL_X1 PHY_226 ();
 AOI221_X1 _05714_ (.A(_01476_),
    .B1(net111),
    .B2(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[15][0] ),
    .C1(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[17][0] ),
    .C2(net81),
    .ZN(_01479_));
 NAND4_X1 _05715_ (.A1(_01463_),
    .A2(_01468_),
    .A3(_01474_),
    .A4(_01479_),
    .ZN(_01480_));
 TAPCELL_X1 PHY_225 ();
 AOI22_X1 _05717_ (.A1(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[24][0] ),
    .A2(_01059_),
    .B1(_01007_),
    .B2(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[13][0] ),
    .ZN(_01482_));
 TAPCELL_X1 PHY_224 ();
 TAPCELL_X1 PHY_223 ();
 TAPCELL_X1 PHY_222 ();
 AOI22_X1 _05721_ (.A1(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[28][0] ),
    .A2(_01032_),
    .B1(net88),
    .B2(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[14][0] ),
    .ZN(_01486_));
 AOI22_X1 _05722_ (.A1(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[27][0] ),
    .A2(net186),
    .B1(net244),
    .B2(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[20][0] ),
    .ZN(_01487_));
 AOI22_X2 _05723_ (.A1(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[16][0] ),
    .A2(net121),
    .B1(net89),
    .B2(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[10][0] ),
    .ZN(_01488_));
 NAND4_X2 _05724_ (.A1(_01482_),
    .A2(_01486_),
    .A3(_01487_),
    .A4(_01488_),
    .ZN(_01489_));
 TAPCELL_X1 PHY_221 ();
 AOI22_X1 _05726_ (.A1(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[5][0] ),
    .A2(net135),
    .B1(_01149_),
    .B2(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[31][0] ),
    .ZN(_01491_));
 AOI22_X1 _05727_ (.A1(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[1][0] ),
    .A2(_00975_),
    .B1(net200),
    .B2(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[19][0] ),
    .ZN(_01492_));
 TAPCELL_X1 PHY_220 ();
 TAPCELL_X1 PHY_219 ();
 TAPCELL_X1 PHY_218 ();
 TAPCELL_X1 PHY_217 ();
 AOI22_X1 _05732_ (.A1(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[29][0] ),
    .A2(_01050_),
    .B1(net228),
    .B2(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[22][0] ),
    .ZN(_01497_));
 TAPCELL_X1 PHY_216 ();
 AOI22_X2 _05734_ (.A1(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[3][0] ),
    .A2(net63),
    .B1(net231),
    .B2(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[11][0] ),
    .ZN(_01499_));
 NAND4_X2 _05735_ (.A1(_01491_),
    .A2(_01492_),
    .A3(_01497_),
    .A4(_01499_),
    .ZN(_01500_));
 NOR3_X2 _05736_ (.A1(_01480_),
    .A2(_01489_),
    .A3(_01500_),
    .ZN(_01501_));
 NOR2_X4 _05737_ (.A1(_00922_),
    .A2(_01407_),
    .ZN(_01502_));
 OAI21_X1 _05738_ (.A(_01502_),
    .B1(net130),
    .B2(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[0][0] ),
    .ZN(_01503_));
 TAPCELL_X1 PHY_215 ();
 AOI22_X1 _05740_ (.A1(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[22][0] ),
    .A2(net224),
    .B1(net219),
    .B2(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[9][0] ),
    .ZN(_01505_));
 AOI22_X1 _05741_ (.A1(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[10][0] ),
    .A2(net90),
    .B1(net241),
    .B2(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[2][0] ),
    .ZN(_01506_));
 AOI22_X1 _05742_ (.A1(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[16][0] ),
    .A2(net117),
    .B1(net170),
    .B2(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[26][0] ),
    .ZN(_01507_));
 AOI22_X2 _05743_ (.A1(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[29][0] ),
    .A2(net142),
    .B1(net269),
    .B2(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[12][0] ),
    .ZN(_01508_));
 NAND4_X2 _05744_ (.A1(_01505_),
    .A2(_01506_),
    .A3(_01507_),
    .A4(_01508_),
    .ZN(_01509_));
 TAPCELL_X1 PHY_214 ();
 AOI22_X1 _05746_ (.A1(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[28][0] ),
    .A2(net77),
    .B1(net68),
    .B2(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[7][0] ),
    .ZN(_01511_));
 TAPCELL_X1 PHY_213 ();
 AOI22_X1 _05748_ (.A1(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[5][0] ),
    .A2(net132),
    .B1(net234),
    .B2(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[11][0] ),
    .ZN(_01513_));
 AOI22_X1 _05749_ (.A1(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[14][0] ),
    .A2(net85),
    .B1(net194),
    .B2(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[19][0] ),
    .ZN(_01514_));
 TAPCELL_X1 PHY_212 ();
 AOI21_X1 _05751_ (.A(net113),
    .B1(net163),
    .B2(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[6][0] ),
    .ZN(_01516_));
 NAND4_X1 _05752_ (.A1(_01511_),
    .A2(_01513_),
    .A3(_01514_),
    .A4(_01516_),
    .ZN(_01517_));
 AOI22_X1 _05753_ (.A1(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[4][0] ),
    .A2(net124),
    .B1(net265),
    .B2(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[18][0] ),
    .ZN(_01518_));
 TAPCELL_X1 PHY_211 ();
 TAPCELL_X1 PHY_210 ();
 AOI22_X1 _05756_ (.A1(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[27][0] ),
    .A2(net190),
    .B1(net74),
    .B2(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[24][0] ),
    .ZN(_01521_));
 TAPCELL_X1 PHY_209 ();
 TAPCELL_X1 PHY_208 ();
 AOI22_X1 _05759_ (.A1(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[31][0] ),
    .A2(net95),
    .B1(net256),
    .B2(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[1][0] ),
    .ZN(_01524_));
 TAPCELL_X1 PHY_207 ();
 AOI22_X1 _05761_ (.A1(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[8][0] ),
    .A2(net179),
    .B1(net209),
    .B2(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[30][0] ),
    .ZN(_01526_));
 NAND4_X1 _05762_ (.A1(_01518_),
    .A2(_01521_),
    .A3(_01524_),
    .A4(_01526_),
    .ZN(_01527_));
 AOI22_X1 _05763_ (.A1(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[17][0] ),
    .A2(net80),
    .B1(net64),
    .B2(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[3][0] ),
    .ZN(_01528_));
 TAPCELL_X1 PHY_206 ();
 TAPCELL_X1 PHY_205 ();
 AOI22_X1 _05766_ (.A1(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[25][0] ),
    .A2(net153),
    .B1(net251),
    .B2(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[20][0] ),
    .ZN(_01531_));
 TAPCELL_X1 PHY_204 ();
 AOI22_X1 _05768_ (.A1(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[15][0] ),
    .A2(net107),
    .B1(net82),
    .B2(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[21][0] ),
    .ZN(_01533_));
 TAPCELL_X1 PHY_203 ();
 TAPCELL_X1 PHY_202 ();
 AOI22_X1 _05771_ (.A1(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[23][0] ),
    .A2(net101),
    .B1(net204),
    .B2(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[13][0] ),
    .ZN(_01536_));
 NAND4_X1 _05772_ (.A1(_01528_),
    .A2(_01531_),
    .A3(_01533_),
    .A4(_01536_),
    .ZN(_01537_));
 NOR4_X2 _05773_ (.A1(_01509_),
    .A2(_01517_),
    .A3(_01527_),
    .A4(_01537_),
    .ZN(_01538_));
 NOR3_X4 _05774_ (.A1(net4),
    .A2(net5),
    .A3(_00921_),
    .ZN(_01539_));
 TAPCELL_X1 PHY_201 ();
 OAI21_X1 _05776_ (.A(_01539_),
    .B1(net130),
    .B2(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[0][0] ),
    .ZN(_01541_));
 OAI22_X1 _05777_ (.A1(_01501_),
    .A2(_01503_),
    .B1(_01538_),
    .B2(_01541_),
    .ZN(_01542_));
 TAPCELL_X1 PHY_200 ();
 AOI22_X1 _05779_ (.A1(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[25][0] ),
    .A2(net147),
    .B1(net229),
    .B2(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[11][0] ),
    .ZN(_01544_));
 TAPCELL_X1 PHY_199 ();
 AOI22_X1 _05781_ (.A1(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[20][0] ),
    .A2(net246),
    .B1(net227),
    .B2(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[22][0] ),
    .ZN(_01546_));
 TAPCELL_X1 PHY_198 ();
 TAPCELL_X1 PHY_197 ();
 TAPCELL_X1 PHY_196 ();
 TAPCELL_X1 PHY_195 ();
 AOI22_X2 _05786_ (.A1(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[16][0] ),
    .A2(net120),
    .B1(net185),
    .B2(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[8][0] ),
    .ZN(_01551_));
 AOI22_X2 _05787_ (.A1(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[6][0] ),
    .A2(net157),
    .B1(net93),
    .B2(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[31][0] ),
    .ZN(_01552_));
 NAND4_X2 _05788_ (.A1(_01544_),
    .A2(_01546_),
    .A3(_01551_),
    .A4(_01552_),
    .ZN(_01553_));
 AOI22_X2 _05789_ (.A1(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[18][0] ),
    .A2(_00964_),
    .B1(net199),
    .B2(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[19][0] ),
    .ZN(_01554_));
 TAPCELL_X1 PHY_194 ();
 TAPCELL_X1 PHY_193 ();
 AOI22_X2 _05792_ (.A1(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[2][0] ),
    .A2(net238),
    .B1(net203),
    .B2(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[13][0] ),
    .ZN(_01557_));
 TAPCELL_X1 PHY_192 ();
 AOI22_X2 _05794_ (.A1(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[15][0] ),
    .A2(net110),
    .B1(net273),
    .B2(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[12][0] ),
    .ZN(_01559_));
 AOI21_X2 _05795_ (.A(net115),
    .B1(_01102_),
    .B2(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[3][0] ),
    .ZN(_01560_));
 NAND4_X4 _05796_ (.A1(_01554_),
    .A2(_01557_),
    .A3(_01559_),
    .A4(_01560_),
    .ZN(_01561_));
 TAPCELL_X1 PHY_191 ();
 AOI22_X1 _05798_ (.A1(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[28][0] ),
    .A2(net76),
    .B1(net83),
    .B2(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[21][0] ),
    .ZN(_01563_));
 TAPCELL_X1 PHY_190 ();
 AOI22_X1 _05800_ (.A1(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[27][0] ),
    .A2(net188),
    .B1(net102),
    .B2(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[23][0] ),
    .ZN(_01565_));
 TAPCELL_X1 PHY_189 ();
 TAPCELL_X1 PHY_188 ();
 AOI22_X1 _05803_ (.A1(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[17][0] ),
    .A2(net79),
    .B1(net218),
    .B2(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[9][0] ),
    .ZN(_01568_));
 TAPCELL_X1 PHY_187 ();
 TAPCELL_X1 PHY_186 ();
 AOI22_X2 _05806_ (.A1(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[29][0] ),
    .A2(net141),
    .B1(net213),
    .B2(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[30][0] ),
    .ZN(_01571_));
 NAND4_X2 _05807_ (.A1(_01563_),
    .A2(_01565_),
    .A3(_01568_),
    .A4(_01571_),
    .ZN(_01572_));
 TAPCELL_X1 PHY_185 ();
 AOI22_X1 _05809_ (.A1(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[7][0] ),
    .A2(net69),
    .B1(net127),
    .B2(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[4][0] ),
    .ZN(_01574_));
 TAPCELL_X1 PHY_184 ();
 AOI22_X1 _05811_ (.A1(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[5][0] ),
    .A2(net133),
    .B1(_01059_),
    .B2(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[24][0] ),
    .ZN(_01576_));
 TAPCELL_X1 PHY_183 ();
 AOI22_X1 _05813_ (.A1(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[14][0] ),
    .A2(net88),
    .B1(net261),
    .B2(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[1][0] ),
    .ZN(_01578_));
 TAPCELL_X1 PHY_182 ();
 AOI22_X2 _05815_ (.A1(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[26][0] ),
    .A2(net166),
    .B1(_00956_),
    .B2(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[10][0] ),
    .ZN(_01580_));
 NAND4_X2 _05816_ (.A1(_01574_),
    .A2(_01576_),
    .A3(_01578_),
    .A4(_01580_),
    .ZN(_01581_));
 NOR4_X4 _05817_ (.A1(_01553_),
    .A2(_01561_),
    .A3(_01572_),
    .A4(_01581_),
    .ZN(_01582_));
 NOR2_X4 _05818_ (.A1(_01163_),
    .A2(_01349_),
    .ZN(_01583_));
 OAI21_X2 _05819_ (.A(_01583_),
    .B1(net130),
    .B2(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[0][0] ),
    .ZN(_01584_));
 TAPCELL_X1 PHY_181 ();
 AOI22_X1 _05821_ (.A1(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[28][0] ),
    .A2(net76),
    .B1(net165),
    .B2(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[6][0] ),
    .ZN(_01586_));
 TAPCELL_X1 PHY_180 ();
 TAPCELL_X1 PHY_179 ();
 AOI22_X1 _05824_ (.A1(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[23][0] ),
    .A2(net97),
    .B1(net110),
    .B2(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[15][0] ),
    .ZN(_01589_));
 TAPCELL_X1 PHY_178 ();
 AOI22_X1 _05826_ (.A1(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[25][0] ),
    .A2(net147),
    .B1(net127),
    .B2(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[4][0] ),
    .ZN(_01591_));
 AOI22_X1 _05827_ (.A1(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[17][0] ),
    .A2(net81),
    .B1(net122),
    .B2(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[16][0] ),
    .ZN(_01592_));
 NAND4_X1 _05828_ (.A1(_01586_),
    .A2(_01589_),
    .A3(_01591_),
    .A4(_01592_),
    .ZN(_01593_));
 TAPCELL_X1 PHY_177 ();
 AOI22_X1 _05830_ (.A1(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[29][0] ),
    .A2(net141),
    .B1(_01059_),
    .B2(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[24][0] ),
    .ZN(_01595_));
 AOI22_X1 _05831_ (.A1(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[27][0] ),
    .A2(net187),
    .B1(net63),
    .B2(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[3][0] ),
    .ZN(_01596_));
 NOR4_X4 _05832_ (.A1(net8),
    .A2(_00953_),
    .A3(net10),
    .A4(_00946_),
    .ZN(_01597_));
 MUX2_X1 _05833_ (.A(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[5][0] ),
    .B(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[21][0] ),
    .S(net1),
    .Z(_01598_));
 TAPCELL_X1 PHY_176 ();
 AOI221_X1 _05835_ (.A(net115),
    .B1(_01597_),
    .B2(_01598_),
    .C1(net203),
    .C2(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[13][0] ),
    .ZN(_01600_));
 NAND3_X1 _05836_ (.A1(_01595_),
    .A2(_01596_),
    .A3(_01600_),
    .ZN(_01601_));
 TAPCELL_X1 PHY_175 ();
 TAPCELL_X1 PHY_174 ();
 AOI22_X1 _05839_ (.A1(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[2][0] ),
    .A2(net239),
    .B1(net202),
    .B2(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[19][0] ),
    .ZN(_01604_));
 TAPCELL_X1 PHY_173 ();
 AOI22_X1 _05841_ (.A1(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[26][0] ),
    .A2(net166),
    .B1(_00964_),
    .B2(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[18][0] ),
    .ZN(_01606_));
 TAPCELL_X1 PHY_172 ();
 AOI22_X1 _05843_ (.A1(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[8][0] ),
    .A2(net177),
    .B1(net70),
    .B2(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[7][0] ),
    .ZN(_01608_));
 AOI22_X2 _05844_ (.A1(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[10][0] ),
    .A2(net89),
    .B1(net261),
    .B2(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[1][0] ),
    .ZN(_01609_));
 NAND4_X2 _05845_ (.A1(_01604_),
    .A2(_01606_),
    .A3(_01608_),
    .A4(_01609_),
    .ZN(_01610_));
 TAPCELL_X1 PHY_171 ();
 TAPCELL_X1 PHY_170 ();
 AOI22_X1 _05848_ (.A1(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[31][0] ),
    .A2(net94),
    .B1(net230),
    .B2(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[11][0] ),
    .ZN(_01613_));
 TAPCELL_X1 PHY_169 ();
 TAPCELL_X1 PHY_168 ();
 AOI22_X1 _05851_ (.A1(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[14][0] ),
    .A2(net88),
    .B1(net246),
    .B2(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[20][0] ),
    .ZN(_01616_));
 AOI22_X1 _05852_ (.A1(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[12][0] ),
    .A2(net273),
    .B1(net218),
    .B2(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[9][0] ),
    .ZN(_01617_));
 TAPCELL_X1 PHY_167 ();
 TAPCELL_X1 PHY_166 ();
 AOI22_X2 _05855_ (.A1(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[22][0] ),
    .A2(net227),
    .B1(net214),
    .B2(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[30][0] ),
    .ZN(_01620_));
 NAND4_X2 _05856_ (.A1(_01613_),
    .A2(_01616_),
    .A3(_01617_),
    .A4(_01620_),
    .ZN(_01621_));
 NOR4_X2 _05857_ (.A1(_01593_),
    .A2(_01601_),
    .A3(_01610_),
    .A4(_01621_),
    .ZN(_01622_));
 NOR3_X4 _05858_ (.A1(net4),
    .A2(net5),
    .A3(_01407_),
    .ZN(_01623_));
 TAPCELL_X1 PHY_165 ();
 OAI21_X1 _05860_ (.A(_01623_),
    .B1(net130),
    .B2(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[0][0] ),
    .ZN(_01625_));
 OAI22_X4 _05861_ (.A1(_01582_),
    .A2(_01584_),
    .B1(_01622_),
    .B2(_01625_),
    .ZN(_01626_));
 TAPCELL_X1 PHY_164 ();
 TAPCELL_X1 PHY_163 ();
 AOI22_X1 _05864_ (.A1(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[18][0] ),
    .A2(_00964_),
    .B1(net262),
    .B2(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[1][0] ),
    .ZN(_01629_));
 TAPCELL_X1 PHY_162 ();
 AOI22_X1 _05866_ (.A1(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[27][0] ),
    .A2(net186),
    .B1(net200),
    .B2(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[19][0] ),
    .ZN(_01631_));
 TAPCELL_X1 PHY_161 ();
 AOI22_X1 _05868_ (.A1(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[15][0] ),
    .A2(net111),
    .B1(net216),
    .B2(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[30][0] ),
    .ZN(_01633_));
 TAPCELL_X1 PHY_160 ();
 AOI22_X2 _05870_ (.A1(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[31][0] ),
    .A2(net94),
    .B1(net129),
    .B2(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[4][0] ),
    .ZN(_01635_));
 NAND4_X2 _05871_ (.A1(_01629_),
    .A2(_01631_),
    .A3(_01633_),
    .A4(_01635_),
    .ZN(_01636_));
 AOI22_X1 _05872_ (.A1(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[16][0] ),
    .A2(net121),
    .B1(net165),
    .B2(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[6][0] ),
    .ZN(_01637_));
 TAPCELL_X1 PHY_159 ();
 AOI22_X1 _05874_ (.A1(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[28][0] ),
    .A2(_01032_),
    .B1(net73),
    .B2(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[24][0] ),
    .ZN(_01639_));
 AOI22_X1 _05875_ (.A1(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[17][0] ),
    .A2(net81),
    .B1(_00986_),
    .B2(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[20][0] ),
    .ZN(_01640_));
 NOR2_X1 _05876_ (.A1(net7),
    .A2(net9),
    .ZN(_01641_));
 NAND2_X1 _05877_ (.A1(net10),
    .A2(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[26][0] ),
    .ZN(_01642_));
 OAI22_X1 _05878_ (.A1(net10),
    .A2(_00948_),
    .B1(_01642_),
    .B2(_00960_),
    .ZN(_01643_));
 AOI22_X1 _05879_ (.A1(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[21][0] ),
    .A2(_00981_),
    .B1(_01641_),
    .B2(_01643_),
    .ZN(_01644_));
 NAND4_X1 _05880_ (.A1(_01637_),
    .A2(_01639_),
    .A3(_01640_),
    .A4(_01644_),
    .ZN(_01645_));
 MUX2_X1 _05881_ (.A(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[5][0] ),
    .B(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[7][0] ),
    .S(net8),
    .Z(_01646_));
 AOI22_X1 _05882_ (.A1(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[23][0] ),
    .A2(_00926_),
    .B1(_01646_),
    .B2(_00911_),
    .ZN(_01647_));
 OR2_X1 _05883_ (.A1(_00980_),
    .A2(_01647_),
    .ZN(_01648_));
 AOI22_X1 _05884_ (.A1(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[25][0] ),
    .A2(net148),
    .B1(net203),
    .B2(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[13][0] ),
    .ZN(_01649_));
 AOI22_X1 _05885_ (.A1(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[12][0] ),
    .A2(_00950_),
    .B1(net218),
    .B2(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[9][0] ),
    .ZN(_01650_));
 NAND3_X1 _05886_ (.A1(_01648_),
    .A2(_01649_),
    .A3(_01650_),
    .ZN(_01651_));
 AOI22_X1 _05887_ (.A1(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[29][0] ),
    .A2(net141),
    .B1(net230),
    .B2(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[11][0] ),
    .ZN(_01652_));
 TAPCELL_X1 PHY_158 ();
 TAPCELL_X1 PHY_157 ();
 AOI22_X1 _05890_ (.A1(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[3][0] ),
    .A2(net63),
    .B1(net88),
    .B2(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[14][0] ),
    .ZN(_01655_));
 TAPCELL_X1 PHY_156 ();
 AOI22_X1 _05892_ (.A1(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[10][0] ),
    .A2(net89),
    .B1(net239),
    .B2(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[2][0] ),
    .ZN(_01657_));
 TAPCELL_X1 PHY_155 ();
 AOI22_X2 _05894_ (.A1(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[8][0] ),
    .A2(net177),
    .B1(net227),
    .B2(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[22][0] ),
    .ZN(_01659_));
 NAND4_X2 _05895_ (.A1(_01652_),
    .A2(_01655_),
    .A3(_01657_),
    .A4(_01659_),
    .ZN(_01660_));
 NOR4_X2 _05896_ (.A1(_01636_),
    .A2(_01645_),
    .A3(_01651_),
    .A4(_01660_),
    .ZN(_01661_));
 NOR3_X4 _05897_ (.A1(net4),
    .A2(net5),
    .A3(_01349_),
    .ZN(_01662_));
 OAI21_X1 _05898_ (.A(_01662_),
    .B1(net130),
    .B2(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[0][0] ),
    .ZN(_01663_));
 TAPCELL_X1 PHY_154 ();
 TAPCELL_X1 PHY_153 ();
 AOI22_X1 _05901_ (.A1(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[4][0] ),
    .A2(net123),
    .B1(net217),
    .B2(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[9][0] ),
    .ZN(_01666_));
 AOI22_X1 _05902_ (.A1(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[29][0] ),
    .A2(net144),
    .B1(net203),
    .B2(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[13][0] ),
    .ZN(_01667_));
 TAPCELL_X1 PHY_152 ();
 AOI22_X1 _05904_ (.A1(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[8][0] ),
    .A2(net178),
    .B1(net175),
    .B2(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[26][0] ),
    .ZN(_01669_));
 AOI22_X1 _05905_ (.A1(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[18][0] ),
    .A2(net263),
    .B1(net236),
    .B2(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[11][0] ),
    .ZN(_01670_));
 NAND4_X1 _05906_ (.A1(_01666_),
    .A2(_01667_),
    .A3(_01669_),
    .A4(_01670_),
    .ZN(_01671_));
 TAPCELL_X1 PHY_151 ();
 AOI22_X1 _05908_ (.A1(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[25][0] ),
    .A2(net152),
    .B1(net196),
    .B2(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[19][0] ),
    .ZN(_01673_));
 AOI22_X1 _05909_ (.A1(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[3][0] ),
    .A2(net64),
    .B1(net260),
    .B2(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[1][0] ),
    .ZN(_01674_));
 TAPCELL_X1 PHY_150 ();
 AOI22_X1 _05911_ (.A1(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[14][0] ),
    .A2(net87),
    .B1(net83),
    .B2(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[21][0] ),
    .ZN(_01676_));
 TAPCELL_X1 PHY_149 ();
 AOI21_X1 _05913_ (.A(net114),
    .B1(net77),
    .B2(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[28][0] ),
    .ZN(_01678_));
 NAND4_X1 _05914_ (.A1(_01673_),
    .A2(_01674_),
    .A3(_01676_),
    .A4(_01678_),
    .ZN(_01679_));
 INV_X1 _05915_ (.A(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[6][0] ),
    .ZN(_01680_));
 NAND4_X4 _05916_ (.A1(_00911_),
    .A2(net8),
    .A3(net9),
    .A4(_00937_),
    .ZN(_01681_));
 INV_X1 _05917_ (.A(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[30][0] ),
    .ZN(_01682_));
 OAI22_X1 _05918_ (.A1(_01680_),
    .A2(_01681_),
    .B1(_01204_),
    .B2(_01682_),
    .ZN(_01683_));
 TAPCELL_X1 PHY_148 ();
 AOI221_X1 _05920_ (.A(_01683_),
    .B1(net242),
    .B2(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[2][0] ),
    .C1(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[10][0] ),
    .C2(net91),
    .ZN(_01685_));
 INV_X1 _05921_ (.A(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[23][0] ),
    .ZN(_01686_));
 INV_X1 _05922_ (.A(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[15][0] ),
    .ZN(_01687_));
 OAI22_X1 _05923_ (.A1(_01686_),
    .A2(_01417_),
    .B1(_01029_),
    .B2(_01687_),
    .ZN(_01688_));
 AOI221_X1 _05924_ (.A(_01688_),
    .B1(net80),
    .B2(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[17][0] ),
    .C1(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[31][0] ),
    .C2(net95),
    .ZN(_01689_));
 INV_X1 _05925_ (.A(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[12][0] ),
    .ZN(_01690_));
 NAND4_X4 _05926_ (.A1(net1),
    .A2(_00978_),
    .A3(net9),
    .A4(_00937_),
    .ZN(_01691_));
 INV_X1 _05927_ (.A(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[20][0] ),
    .ZN(_01692_));
 OAI22_X1 _05928_ (.A1(_01690_),
    .A2(_01426_),
    .B1(_01691_),
    .B2(_01692_),
    .ZN(_01693_));
 AOI221_X1 _05929_ (.A(_01693_),
    .B1(_01076_),
    .B2(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[7][0] ),
    .C1(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[24][0] ),
    .C2(net72),
    .ZN(_01694_));
 AOI22_X1 _05930_ (.A1(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[27][0] ),
    .A2(net192),
    .B1(net226),
    .B2(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[22][0] ),
    .ZN(_01695_));
 AOI22_X1 _05931_ (.A1(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[16][0] ),
    .A2(net120),
    .B1(net134),
    .B2(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[5][0] ),
    .ZN(_01696_));
 AND2_X1 _05932_ (.A1(_01695_),
    .A2(_01696_),
    .ZN(_01697_));
 NAND4_X1 _05933_ (.A1(_01685_),
    .A2(_01689_),
    .A3(_01694_),
    .A4(_01697_),
    .ZN(_01698_));
 NOR3_X1 _05934_ (.A1(_01671_),
    .A2(_01679_),
    .A3(_01698_),
    .ZN(_01699_));
 NOR2_X4 _05935_ (.A1(_00921_),
    .A2(_01163_),
    .ZN(_01700_));
 TAPCELL_X1 PHY_147 ();
 OAI21_X1 _05937_ (.A(_01700_),
    .B1(net130),
    .B2(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[0][0] ),
    .ZN(_01702_));
 OAI22_X1 _05938_ (.A1(_01661_),
    .A2(_01663_),
    .B1(_01699_),
    .B2(_01702_),
    .ZN(_01703_));
 AOI22_X2 _05939_ (.A1(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[8][0] ),
    .A2(net176),
    .B1(net264),
    .B2(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[18][0] ),
    .ZN(_01704_));
 AOI22_X2 _05940_ (.A1(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[28][0] ),
    .A2(_01032_),
    .B1(net135),
    .B2(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[5][0] ),
    .ZN(_01705_));
 AOI22_X2 _05941_ (.A1(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[1][0] ),
    .A2(net253),
    .B1(_00989_),
    .B2(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[2][0] ),
    .ZN(_01706_));
 AOI22_X2 _05942_ (.A1(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[17][0] ),
    .A2(net81),
    .B1(net186),
    .B2(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[27][0] ),
    .ZN(_01707_));
 NAND4_X4 _05943_ (.A1(_01704_),
    .A2(_01705_),
    .A3(_01706_),
    .A4(_01707_),
    .ZN(_01708_));
 AOI22_X1 _05944_ (.A1(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[23][0] ),
    .A2(net99),
    .B1(_00999_),
    .B2(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[9][0] ),
    .ZN(_01709_));
 AOI22_X1 _05945_ (.A1(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[12][0] ),
    .A2(net272),
    .B1(net244),
    .B2(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[20][0] ),
    .ZN(_01710_));
 TAPCELL_X1 PHY_146 ();
 AOI21_X1 _05947_ (.A(net115),
    .B1(net228),
    .B2(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[22][0] ),
    .ZN(_01712_));
 AOI22_X2 _05948_ (.A1(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[7][0] ),
    .A2(net70),
    .B1(net237),
    .B2(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[11][0] ),
    .ZN(_01713_));
 NAND4_X2 _05949_ (.A1(_01709_),
    .A2(_01710_),
    .A3(_01712_),
    .A4(_01713_),
    .ZN(_01714_));
 AOI22_X1 _05950_ (.A1(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[31][0] ),
    .A2(_01149_),
    .B1(net84),
    .B2(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[21][0] ),
    .ZN(_01715_));
 AOI22_X1 _05951_ (.A1(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[6][0] ),
    .A2(net156),
    .B1(net89),
    .B2(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[10][0] ),
    .ZN(_01716_));
 TAPCELL_X1 PHY_145 ();
 AOI22_X1 _05953_ (.A1(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[29][0] ),
    .A2(net146),
    .B1(net73),
    .B2(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[24][0] ),
    .ZN(_01718_));
 TAPCELL_X1 PHY_144 ();
 TAPCELL_X1 PHY_143 ();
 AOI22_X2 _05956_ (.A1(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[15][0] ),
    .A2(net112),
    .B1(net171),
    .B2(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[26][0] ),
    .ZN(_01721_));
 NAND4_X2 _05957_ (.A1(_01715_),
    .A2(_01716_),
    .A3(_01718_),
    .A4(_01721_),
    .ZN(_01722_));
 AOI22_X1 _05958_ (.A1(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[4][0] ),
    .A2(net128),
    .B1(net206),
    .B2(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[13][0] ),
    .ZN(_01723_));
 TAPCELL_X1 PHY_142 ();
 AOI22_X1 _05960_ (.A1(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[3][0] ),
    .A2(net63),
    .B1(_00971_),
    .B2(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[14][0] ),
    .ZN(_01725_));
 TAPCELL_X1 PHY_141 ();
 AOI22_X1 _05962_ (.A1(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[16][0] ),
    .A2(net121),
    .B1(net150),
    .B2(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[25][0] ),
    .ZN(_01727_));
 AOI22_X2 _05963_ (.A1(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[30][0] ),
    .A2(net215),
    .B1(net201),
    .B2(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[19][0] ),
    .ZN(_01728_));
 NAND4_X2 _05964_ (.A1(_01723_),
    .A2(_01725_),
    .A3(_01727_),
    .A4(_01728_),
    .ZN(_01729_));
 NOR4_X4 _05965_ (.A1(_01708_),
    .A2(_01714_),
    .A3(_01722_),
    .A4(_01729_),
    .ZN(_01730_));
 NOR3_X4 _05966_ (.A1(net2),
    .A2(net3),
    .A3(_00922_),
    .ZN(_01731_));
 TAPCELL_X1 PHY_140 ();
 OAI21_X1 _05968_ (.A(_01731_),
    .B1(net130),
    .B2(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[0][0] ),
    .ZN(_01733_));
 AOI22_X1 _05969_ (.A1(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[31][0] ),
    .A2(net96),
    .B1(net83),
    .B2(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[21][0] ),
    .ZN(_01734_));
 AOI22_X1 _05970_ (.A1(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[17][0] ),
    .A2(net78),
    .B1(_00950_),
    .B2(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[12][0] ),
    .ZN(_01735_));
 AOI22_X1 _05971_ (.A1(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[2][0] ),
    .A2(net241),
    .B1(net235),
    .B2(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[11][0] ),
    .ZN(_01736_));
 AOI22_X1 _05972_ (.A1(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[14][0] ),
    .A2(net87),
    .B1(net205),
    .B2(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[13][0] ),
    .ZN(_01737_));
 NAND4_X1 _05973_ (.A1(_01734_),
    .A2(_01735_),
    .A3(_01736_),
    .A4(_01737_),
    .ZN(_01738_));
 TAPCELL_X1 PHY_139 ();
 AOI22_X1 _05975_ (.A1(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[3][0] ),
    .A2(net65),
    .B1(net72),
    .B2(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[24][0] ),
    .ZN(_01740_));
 TAPCELL_X1 PHY_138 ();
 AOI22_X1 _05977_ (.A1(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[5][0] ),
    .A2(net138),
    .B1(net68),
    .B2(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[7][0] ),
    .ZN(_01742_));
 TAPCELL_X1 PHY_137 ();
 AOI22_X1 _05979_ (.A1(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[9][0] ),
    .A2(net221),
    .B1(_01009_),
    .B2(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[19][0] ),
    .ZN(_01744_));
 TAPCELL_X1 PHY_136 ();
 TAPCELL_X1 PHY_135 ();
 AOI21_X1 _05982_ (.A(net114),
    .B1(net75),
    .B2(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[28][0] ),
    .ZN(_01747_));
 NAND4_X1 _05983_ (.A1(_01740_),
    .A2(_01742_),
    .A3(_01744_),
    .A4(_01747_),
    .ZN(_01748_));
 TAPCELL_X1 PHY_134 ();
 AOI22_X1 _05985_ (.A1(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[15][0] ),
    .A2(net108),
    .B1(net164),
    .B2(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[6][0] ),
    .ZN(_01750_));
 AOI22_X1 _05986_ (.A1(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[27][0] ),
    .A2(net192),
    .B1(_01034_),
    .B2(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[8][0] ),
    .ZN(_01751_));
 TAPCELL_X1 PHY_133 ();
 AOI22_X1 _05988_ (.A1(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[1][0] ),
    .A2(_00975_),
    .B1(net225),
    .B2(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[22][0] ),
    .ZN(_01753_));
 AOI22_X1 _05989_ (.A1(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[16][0] ),
    .A2(_01097_),
    .B1(net211),
    .B2(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[30][0] ),
    .ZN(_01754_));
 NAND4_X1 _05990_ (.A1(_01750_),
    .A2(_01751_),
    .A3(_01753_),
    .A4(_01754_),
    .ZN(_01755_));
 TAPCELL_X1 PHY_132 ();
 AOI22_X1 _05992_ (.A1(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[29][0] ),
    .A2(net143),
    .B1(net249),
    .B2(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[20][0] ),
    .ZN(_01757_));
 TAPCELL_X1 PHY_131 ();
 AOI22_X1 _05994_ (.A1(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[4][0] ),
    .A2(net125),
    .B1(net265),
    .B2(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[18][0] ),
    .ZN(_01759_));
 AOI22_X1 _05995_ (.A1(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[23][0] ),
    .A2(net105),
    .B1(net91),
    .B2(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[10][0] ),
    .ZN(_01760_));
 AOI22_X1 _05996_ (.A1(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[26][0] ),
    .A2(net170),
    .B1(net155),
    .B2(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[25][0] ),
    .ZN(_01761_));
 NAND4_X1 _05997_ (.A1(_01757_),
    .A2(_01759_),
    .A3(_01760_),
    .A4(_01761_),
    .ZN(_01762_));
 NOR4_X1 _05998_ (.A1(_01738_),
    .A2(_01748_),
    .A3(_01755_),
    .A4(_01762_),
    .ZN(_01763_));
 NOR2_X2 _05999_ (.A1(_01163_),
    .A2(_01407_),
    .ZN(_01764_));
 TAPCELL_X1 PHY_130 ();
 OAI21_X1 _06001_ (.A(_01764_),
    .B1(net130),
    .B2(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[0][0] ),
    .ZN(_01766_));
 OAI22_X2 _06002_ (.A1(_01730_),
    .A2(_01733_),
    .B1(_01763_),
    .B2(_01766_),
    .ZN(_01767_));
 NOR4_X2 _06003_ (.A1(_01542_),
    .A2(_01626_),
    .A3(_01703_),
    .A4(_01767_),
    .ZN(_01768_));
 TAPCELL_X1 PHY_129 ();
 TAPCELL_X1 PHY_128 ();
 TAPCELL_X1 PHY_127 ();
 AOI22_X1 _06007_ (.A1(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[26][0] ),
    .A2(net173),
    .B1(net90),
    .B2(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[10][0] ),
    .ZN(_01772_));
 TAPCELL_X1 PHY_126 ();
 TAPCELL_X1 PHY_125 ();
 AOI22_X1 _06010_ (.A1(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[3][0] ),
    .A2(net64),
    .B1(net85),
    .B2(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[14][0] ),
    .ZN(_01775_));
 TAPCELL_X1 PHY_124 ();
 TAPCELL_X1 PHY_123 ();
 AOI22_X1 _06013_ (.A1(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[8][0] ),
    .A2(net179),
    .B1(net250),
    .B2(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[20][0] ),
    .ZN(_01778_));
 TAPCELL_X1 PHY_122 ();
 TAPCELL_X1 PHY_121 ();
 AOI22_X1 _06016_ (.A1(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[27][0] ),
    .A2(net190),
    .B1(net153),
    .B2(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[25][0] ),
    .ZN(_01781_));
 NAND4_X1 _06017_ (.A1(_01772_),
    .A2(_01775_),
    .A3(_01778_),
    .A4(_01781_),
    .ZN(_01782_));
 TAPCELL_X1 PHY_120 ();
 TAPCELL_X1 PHY_119 ();
 AOI22_X1 _06020_ (.A1(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[23][0] ),
    .A2(net100),
    .B1(net116),
    .B2(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[16][0] ),
    .ZN(_01785_));
 TAPCELL_X1 PHY_118 ();
 AOI22_X1 _06022_ (.A1(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[17][0] ),
    .A2(net79),
    .B1(net219),
    .B2(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[9][0] ),
    .ZN(_01787_));
 TAPCELL_X1 PHY_117 ();
 TAPCELL_X1 PHY_116 ();
 AOI22_X1 _06025_ (.A1(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[30][0] ),
    .A2(net209),
    .B1(net204),
    .B2(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[13][0] ),
    .ZN(_01790_));
 TAPCELL_X1 PHY_115 ();
 TAPCELL_X1 PHY_114 ();
 AOI21_X1 _06028_ (.A(net113),
    .B1(net194),
    .B2(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[19][0] ),
    .ZN(_01793_));
 NAND4_X1 _06029_ (.A1(_01785_),
    .A2(_01787_),
    .A3(_01790_),
    .A4(_01793_),
    .ZN(_01794_));
 TAPCELL_X1 PHY_113 ();
 TAPCELL_X1 PHY_112 ();
 AOI22_X1 _06032_ (.A1(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[15][0] ),
    .A2(net107),
    .B1(net93),
    .B2(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[31][0] ),
    .ZN(_01797_));
 TAPCELL_X1 PHY_111 ();
 TAPCELL_X1 PHY_110 ();
 TAPCELL_X1 PHY_109 ();
 AOI22_X1 _06036_ (.A1(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[5][0] ),
    .A2(net131),
    .B1(net82),
    .B2(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[21][0] ),
    .ZN(_01801_));
 TAPCELL_X1 PHY_108 ();
 AOI22_X1 _06038_ (.A1(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[29][0] ),
    .A2(net142),
    .B1(net255),
    .B2(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[1][0] ),
    .ZN(_01803_));
 TAPCELL_X1 PHY_107 ();
 AOI22_X1 _06040_ (.A1(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[7][0] ),
    .A2(net68),
    .B1(net233),
    .B2(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[11][0] ),
    .ZN(_01805_));
 NAND4_X1 _06041_ (.A1(_01797_),
    .A2(_01801_),
    .A3(_01803_),
    .A4(_01805_),
    .ZN(_01806_));
 TAPCELL_X1 PHY_106 ();
 TAPCELL_X1 PHY_105 ();
 AOI22_X1 _06044_ (.A1(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[24][0] ),
    .A2(net71),
    .B1(net240),
    .B2(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[2][0] ),
    .ZN(_01809_));
 TAPCELL_X1 PHY_104 ();
 AOI22_X1 _06046_ (.A1(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[4][0] ),
    .A2(net123),
    .B1(net263),
    .B2(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[18][0] ),
    .ZN(_01811_));
 AOI22_X1 _06047_ (.A1(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[12][0] ),
    .A2(net267),
    .B1(net226),
    .B2(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[22][0] ),
    .ZN(_01812_));
 TAPCELL_X1 PHY_103 ();
 TAPCELL_X1 PHY_102 ();
 AOI22_X2 _06050_ (.A1(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[28][0] ),
    .A2(net76),
    .B1(net162),
    .B2(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[6][0] ),
    .ZN(_01815_));
 NAND4_X2 _06051_ (.A1(_01809_),
    .A2(_01811_),
    .A3(_01812_),
    .A4(_01815_),
    .ZN(_01816_));
 OR4_X2 _06052_ (.A1(_01782_),
    .A2(_01794_),
    .A3(_01806_),
    .A4(_01816_),
    .ZN(_01817_));
 TAPCELL_X1 PHY_101 ();
 OAI21_X1 _06054_ (.A(_01817_),
    .B1(net130),
    .B2(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[0][0] ),
    .ZN(_01819_));
 NOR4_X4 _06055_ (.A1(net2),
    .A2(net3),
    .A3(net4),
    .A4(net5),
    .ZN(_01820_));
 AOI221_X2 _06056_ (.A(_00907_),
    .B1(_01458_),
    .B2(_01768_),
    .C1(_01819_),
    .C2(_01820_),
    .ZN(\rdata_o_n[0] ));
 AOI22_X1 _06057_ (.A1(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[17][1] ),
    .A2(net81),
    .B1(net227),
    .B2(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[22][1] ),
    .ZN(_01821_));
 AOI22_X1 _06058_ (.A1(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[16][1] ),
    .A2(net122),
    .B1(net216),
    .B2(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[30][1] ),
    .ZN(_01822_));
 AOI22_X1 _06059_ (.A1(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[9][1] ),
    .A2(net218),
    .B1(net203),
    .B2(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[13][1] ),
    .ZN(_01823_));
 AOI22_X1 _06060_ (.A1(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[26][1] ),
    .A2(net166),
    .B1(net127),
    .B2(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[4][1] ),
    .ZN(_01824_));
 NAND4_X1 _06061_ (.A1(_01821_),
    .A2(_01822_),
    .A3(_01823_),
    .A4(_01824_),
    .ZN(_01825_));
 AOI22_X1 _06062_ (.A1(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[27][1] ),
    .A2(net187),
    .B1(net147),
    .B2(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[25][1] ),
    .ZN(_01826_));
 AOI22_X1 _06063_ (.A1(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[5][1] ),
    .A2(net133),
    .B1(net261),
    .B2(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[1][1] ),
    .ZN(_01827_));
 TAPCELL_X1 PHY_100 ();
 MUX2_X1 _06065_ (.A(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[12][1] ),
    .B(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[14][1] ),
    .S(net8),
    .Z(_01829_));
 AOI221_X1 _06066_ (.A(net115),
    .B1(net92),
    .B2(_01829_),
    .C1(net230),
    .C2(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[11][1] ),
    .ZN(_01830_));
 NAND3_X1 _06067_ (.A1(_01826_),
    .A2(_01827_),
    .A3(_01830_),
    .ZN(_01831_));
 TAPCELL_X1 PHY_99 ();
 AOI22_X1 _06069_ (.A1(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[15][1] ),
    .A2(net110),
    .B1(_01059_),
    .B2(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[24][1] ),
    .ZN(_01833_));
 AOI22_X1 _06070_ (.A1(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[10][1] ),
    .A2(net89),
    .B1(net202),
    .B2(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[19][1] ),
    .ZN(_01834_));
 TAPCELL_X1 PHY_98 ();
 AOI22_X1 _06072_ (.A1(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[28][1] ),
    .A2(net76),
    .B1(net246),
    .B2(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[20][1] ),
    .ZN(_01836_));
 AOI22_X1 _06073_ (.A1(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[31][1] ),
    .A2(net94),
    .B1(_00964_),
    .B2(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[18][1] ),
    .ZN(_01837_));
 NAND4_X1 _06074_ (.A1(_01833_),
    .A2(_01834_),
    .A3(_01836_),
    .A4(_01837_),
    .ZN(_01838_));
 AOI22_X1 _06075_ (.A1(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[29][1] ),
    .A2(net141),
    .B1(_00981_),
    .B2(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[21][1] ),
    .ZN(_01839_));
 AOI22_X1 _06076_ (.A1(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[23][1] ),
    .A2(net97),
    .B1(net70),
    .B2(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[7][1] ),
    .ZN(_01840_));
 AOI22_X1 _06077_ (.A1(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[8][1] ),
    .A2(net177),
    .B1(net239),
    .B2(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[2][1] ),
    .ZN(_01841_));
 TAPCELL_X1 PHY_97 ();
 AOI22_X2 _06079_ (.A1(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[3][1] ),
    .A2(net63),
    .B1(net159),
    .B2(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[6][1] ),
    .ZN(_01843_));
 NAND4_X2 _06080_ (.A1(_01839_),
    .A2(_01840_),
    .A3(_01841_),
    .A4(_01843_),
    .ZN(_01844_));
 NOR4_X2 _06081_ (.A1(_01825_),
    .A2(_01831_),
    .A3(_01838_),
    .A4(_01844_),
    .ZN(_01845_));
 OAI21_X1 _06082_ (.A(_01623_),
    .B1(net130),
    .B2(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[0][1] ),
    .ZN(_01846_));
 AOI22_X1 _06083_ (.A1(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[3][1] ),
    .A2(net65),
    .B1(_01042_),
    .B2(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[6][1] ),
    .ZN(_01847_));
 TAPCELL_X1 PHY_96 ();
 AOI22_X1 _06085_ (.A1(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[12][1] ),
    .A2(net272),
    .B1(net243),
    .B2(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[2][1] ),
    .ZN(_01849_));
 AOI22_X1 _06086_ (.A1(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[14][1] ),
    .A2(net87),
    .B1(net206),
    .B2(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[13][1] ),
    .ZN(_01850_));
 AOI22_X1 _06087_ (.A1(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[17][1] ),
    .A2(net78),
    .B1(net183),
    .B2(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[8][1] ),
    .ZN(_01851_));
 NAND4_X1 _06088_ (.A1(_01847_),
    .A2(_01849_),
    .A3(_01850_),
    .A4(_01851_),
    .ZN(_01852_));
 TAPCELL_X1 PHY_95 ();
 AOI22_X1 _06090_ (.A1(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[7][1] ),
    .A2(net70),
    .B1(net211),
    .B2(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[30][1] ),
    .ZN(_01854_));
 AOI22_X1 _06091_ (.A1(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[25][1] ),
    .A2(net150),
    .B1(_00999_),
    .B2(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[9][1] ),
    .ZN(_01855_));
 TAPCELL_X1 PHY_94 ();
 AOI21_X1 _06093_ (.A(net115),
    .B1(_01149_),
    .B2(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[31][1] ),
    .ZN(_01857_));
 AOI22_X1 _06094_ (.A1(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[16][1] ),
    .A2(net119),
    .B1(net201),
    .B2(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[19][1] ),
    .ZN(_01858_));
 NAND4_X1 _06095_ (.A1(_01854_),
    .A2(_01855_),
    .A3(_01857_),
    .A4(_01858_),
    .ZN(_01859_));
 AOI22_X1 _06096_ (.A1(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[29][1] ),
    .A2(net146),
    .B1(net253),
    .B2(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[1][1] ),
    .ZN(_01860_));
 AOI22_X1 _06097_ (.A1(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[15][1] ),
    .A2(net109),
    .B1(net264),
    .B2(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[18][1] ),
    .ZN(_01861_));
 AOI22_X1 _06098_ (.A1(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[28][1] ),
    .A2(_01032_),
    .B1(net171),
    .B2(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[26][1] ),
    .ZN(_01862_));
 TAPCELL_X1 PHY_93 ();
 AOI22_X2 _06100_ (.A1(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[23][1] ),
    .A2(net99),
    .B1(net73),
    .B2(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[24][1] ),
    .ZN(_01864_));
 NAND4_X2 _06101_ (.A1(_01860_),
    .A2(_01861_),
    .A3(_01862_),
    .A4(_01864_),
    .ZN(_01865_));
 TAPCELL_X1 PHY_92 ();
 AOI22_X1 _06103_ (.A1(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[20][1] ),
    .A2(net252),
    .B1(net225),
    .B2(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[22][1] ),
    .ZN(_01867_));
 TAPCELL_X1 PHY_91 ();
 AOI22_X1 _06105_ (.A1(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[27][1] ),
    .A2(net192),
    .B1(net139),
    .B2(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[5][1] ),
    .ZN(_01869_));
 TAPCELL_X1 PHY_90 ();
 AOI22_X1 _06107_ (.A1(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[21][1] ),
    .A2(net84),
    .B1(net237),
    .B2(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[11][1] ),
    .ZN(_01871_));
 TAPCELL_X1 PHY_89 ();
 AOI22_X1 _06109_ (.A1(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[4][1] ),
    .A2(net128),
    .B1(net89),
    .B2(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[10][1] ),
    .ZN(_01873_));
 NAND4_X1 _06110_ (.A1(_01867_),
    .A2(_01869_),
    .A3(_01871_),
    .A4(_01873_),
    .ZN(_01874_));
 NOR4_X2 _06111_ (.A1(_01852_),
    .A2(_01859_),
    .A3(_01865_),
    .A4(_01874_),
    .ZN(_01875_));
 OAI21_X1 _06112_ (.A(_01408_),
    .B1(net130),
    .B2(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[0][1] ),
    .ZN(_01876_));
 OAI22_X2 _06113_ (.A1(_01845_),
    .A2(_01846_),
    .B1(_01875_),
    .B2(_01876_),
    .ZN(_01877_));
 AOI22_X1 _06114_ (.A1(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[31][1] ),
    .A2(net95),
    .B1(net234),
    .B2(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[11][1] ),
    .ZN(_01878_));
 AOI22_X1 _06115_ (.A1(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[28][1] ),
    .A2(net77),
    .B1(net82),
    .B2(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[21][1] ),
    .ZN(_01879_));
 AOI22_X1 _06116_ (.A1(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[17][1] ),
    .A2(net80),
    .B1(net132),
    .B2(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[5][1] ),
    .ZN(_01880_));
 AOI22_X1 _06117_ (.A1(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[12][1] ),
    .A2(net269),
    .B1(net85),
    .B2(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[14][1] ),
    .ZN(_01881_));
 NAND4_X1 _06118_ (.A1(_01878_),
    .A2(_01879_),
    .A3(_01880_),
    .A4(_01881_),
    .ZN(_01882_));
 AOI22_X1 _06119_ (.A1(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[8][1] ),
    .A2(net181),
    .B1(net204),
    .B2(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[13][1] ),
    .ZN(_01883_));
 AOI22_X1 _06120_ (.A1(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[6][1] ),
    .A2(net163),
    .B1(net68),
    .B2(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[7][1] ),
    .ZN(_01884_));
 AOI22_X1 _06121_ (.A1(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[29][1] ),
    .A2(net142),
    .B1(net251),
    .B2(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[20][1] ),
    .ZN(_01885_));
 AOI21_X1 _06122_ (.A(net113),
    .B1(net256),
    .B2(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[1][1] ),
    .ZN(_01886_));
 NAND4_X1 _06123_ (.A1(_01883_),
    .A2(_01884_),
    .A3(_01885_),
    .A4(_01886_),
    .ZN(_01887_));
 AOI22_X1 _06124_ (.A1(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[15][1] ),
    .A2(net106),
    .B1(net209),
    .B2(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[30][1] ),
    .ZN(_01888_));
 AOI22_X1 _06125_ (.A1(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[3][1] ),
    .A2(net64),
    .B1(net219),
    .B2(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[9][1] ),
    .ZN(_01889_));
 AOI22_X1 _06126_ (.A1(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[4][1] ),
    .A2(net124),
    .B1(net224),
    .B2(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[22][1] ),
    .ZN(_01890_));
 TAPCELL_X1 PHY_88 ();
 AOI22_X1 _06128_ (.A1(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[25][1] ),
    .A2(net153),
    .B1(net265),
    .B2(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[18][1] ),
    .ZN(_01892_));
 NAND4_X1 _06129_ (.A1(_01888_),
    .A2(_01889_),
    .A3(_01890_),
    .A4(_01892_),
    .ZN(_01893_));
 AOI22_X1 _06130_ (.A1(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[10][1] ),
    .A2(net90),
    .B1(net195),
    .B2(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[19][1] ),
    .ZN(_01894_));
 AOI22_X1 _06131_ (.A1(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[27][1] ),
    .A2(net190),
    .B1(net170),
    .B2(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[26][1] ),
    .ZN(_01895_));
 TAPCELL_X1 PHY_87 ();
 AOI22_X1 _06133_ (.A1(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[23][1] ),
    .A2(net101),
    .B1(net117),
    .B2(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[16][1] ),
    .ZN(_01897_));
 AOI22_X1 _06134_ (.A1(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[24][1] ),
    .A2(net74),
    .B1(net241),
    .B2(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[2][1] ),
    .ZN(_01898_));
 NAND4_X1 _06135_ (.A1(_01894_),
    .A2(_01895_),
    .A3(_01897_),
    .A4(_01898_),
    .ZN(_01899_));
 NOR4_X1 _06136_ (.A1(_01882_),
    .A2(_01887_),
    .A3(_01893_),
    .A4(_01899_),
    .ZN(_01900_));
 OAI21_X1 _06137_ (.A(_01539_),
    .B1(net130),
    .B2(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[0][1] ),
    .ZN(_01901_));
 OAI21_X1 _06138_ (.A(_01406_),
    .B1(_01900_),
    .B2(_01901_),
    .ZN(_01902_));
 AOI22_X1 _06139_ (.A1(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[17][1] ),
    .A2(net81),
    .B1(net246),
    .B2(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[20][1] ),
    .ZN(_01903_));
 AOI221_X1 _06140_ (.A(net115),
    .B1(net261),
    .B2(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[1][1] ),
    .C1(net199),
    .C2(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[19][1] ),
    .ZN(_01904_));
 AOI22_X1 _06141_ (.A1(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[27][1] ),
    .A2(net187),
    .B1(_00964_),
    .B2(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[18][1] ),
    .ZN(_01905_));
 AOI22_X1 _06142_ (.A1(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[16][1] ),
    .A2(net122),
    .B1(net227),
    .B2(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[22][1] ),
    .ZN(_01906_));
 NAND4_X1 _06143_ (.A1(_01903_),
    .A2(_01904_),
    .A3(_01905_),
    .A4(_01906_),
    .ZN(_01907_));
 AOI22_X1 _06144_ (.A1(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[12][1] ),
    .A2(net273),
    .B1(net88),
    .B2(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[14][1] ),
    .ZN(_01908_));
 TAPCELL_X1 PHY_86 ();
 AOI22_X1 _06146_ (.A1(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[25][1] ),
    .A2(net147),
    .B1(net69),
    .B2(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[7][1] ),
    .ZN(_01910_));
 AOI22_X1 _06147_ (.A1(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[5][1] ),
    .A2(net133),
    .B1(net94),
    .B2(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[31][1] ),
    .ZN(_01911_));
 AOI22_X1 _06148_ (.A1(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[23][1] ),
    .A2(net97),
    .B1(_00981_),
    .B2(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[21][1] ),
    .ZN(_01912_));
 NAND4_X1 _06149_ (.A1(_01908_),
    .A2(_01910_),
    .A3(_01911_),
    .A4(_01912_),
    .ZN(_01913_));
 TAPCELL_X1 PHY_85 ();
 AOI22_X1 _06151_ (.A1(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[6][1] ),
    .A2(net157),
    .B1(net218),
    .B2(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[9][1] ),
    .ZN(_01915_));
 AOI22_X1 _06152_ (.A1(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[28][1] ),
    .A2(net76),
    .B1(net238),
    .B2(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[2][1] ),
    .ZN(_01916_));
 AOI22_X1 _06153_ (.A1(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[15][1] ),
    .A2(net110),
    .B1(_00956_),
    .B2(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[10][1] ),
    .ZN(_01917_));
 AOI22_X1 _06154_ (.A1(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[8][1] ),
    .A2(net185),
    .B1(net141),
    .B2(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[29][1] ),
    .ZN(_01918_));
 NAND4_X1 _06155_ (.A1(_01915_),
    .A2(_01916_),
    .A3(_01917_),
    .A4(_01918_),
    .ZN(_01919_));
 TAPCELL_X1 PHY_84 ();
 AOI22_X1 _06157_ (.A1(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[3][1] ),
    .A2(_01102_),
    .B1(net203),
    .B2(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[13][1] ),
    .ZN(_01921_));
 AOI222_X2 _06158_ (.A1(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[26][1] ),
    .A2(net166),
    .B1(_01059_),
    .B2(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[24][1] ),
    .C1(net230),
    .C2(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[11][1] ),
    .ZN(_01922_));
 AOI22_X1 _06159_ (.A1(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[4][1] ),
    .A2(net127),
    .B1(net214),
    .B2(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[30][1] ),
    .ZN(_01923_));
 NAND3_X1 _06160_ (.A1(_01921_),
    .A2(_01922_),
    .A3(_01923_),
    .ZN(_01924_));
 NOR4_X2 _06161_ (.A1(_01907_),
    .A2(_01913_),
    .A3(_01919_),
    .A4(_01924_),
    .ZN(_01925_));
 OAI21_X1 _06162_ (.A(_01583_),
    .B1(net130),
    .B2(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[0][1] ),
    .ZN(_01926_));
 AOI22_X1 _06163_ (.A1(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[16][1] ),
    .A2(net120),
    .B1(net87),
    .B2(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[14][1] ),
    .ZN(_01927_));
 AOI22_X1 _06164_ (.A1(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[8][1] ),
    .A2(net178),
    .B1(net254),
    .B2(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[1][1] ),
    .ZN(_01928_));
 AOI22_X1 _06165_ (.A1(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[23][1] ),
    .A2(net102),
    .B1(net93),
    .B2(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[31][1] ),
    .ZN(_01929_));
 TAPCELL_X1 PHY_83 ();
 AOI22_X2 _06167_ (.A1(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[7][1] ),
    .A2(net69),
    .B1(net245),
    .B2(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[20][1] ),
    .ZN(_01931_));
 NAND4_X2 _06168_ (.A1(_01927_),
    .A2(_01928_),
    .A3(_01929_),
    .A4(_01931_),
    .ZN(_01932_));
 AOI22_X1 _06169_ (.A1(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[15][1] ),
    .A2(net110),
    .B1(net158),
    .B2(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[6][1] ),
    .ZN(_01933_));
 AOI22_X1 _06170_ (.A1(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[4][1] ),
    .A2(net126),
    .B1(net268),
    .B2(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[12][1] ),
    .ZN(_01934_));
 TAPCELL_X1 PHY_82 ();
 AOI22_X1 _06172_ (.A1(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[27][1] ),
    .A2(net188),
    .B1(net144),
    .B2(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[29][1] ),
    .ZN(_01936_));
 AOI21_X1 _06173_ (.A(net114),
    .B1(net66),
    .B2(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[3][1] ),
    .ZN(_01937_));
 NAND4_X1 _06174_ (.A1(_01933_),
    .A2(_01934_),
    .A3(_01936_),
    .A4(_01937_),
    .ZN(_01938_));
 AOI22_X1 _06175_ (.A1(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[26][1] ),
    .A2(net174),
    .B1(net196),
    .B2(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[19][1] ),
    .ZN(_01939_));
 AOI22_X1 _06176_ (.A1(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[10][1] ),
    .A2(_00956_),
    .B1(net263),
    .B2(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[18][1] ),
    .ZN(_01940_));
 TAPCELL_X1 PHY_81 ();
 AOI22_X1 _06178_ (.A1(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[25][1] ),
    .A2(net148),
    .B1(net217),
    .B2(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[9][1] ),
    .ZN(_01942_));
 TAPCELL_X1 PHY_80 ();
 AOI22_X1 _06180_ (.A1(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[24][1] ),
    .A2(net71),
    .B1(net83),
    .B2(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[21][1] ),
    .ZN(_01944_));
 NAND4_X1 _06181_ (.A1(_01939_),
    .A2(_01940_),
    .A3(_01942_),
    .A4(_01944_),
    .ZN(_01945_));
 TAPCELL_X1 PHY_79 ();
 AOI22_X1 _06183_ (.A1(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[28][1] ),
    .A2(net76),
    .B1(net238),
    .B2(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[2][1] ),
    .ZN(_01947_));
 AOI22_X1 _06184_ (.A1(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[11][1] ),
    .A2(net229),
    .B1(net203),
    .B2(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[13][1] ),
    .ZN(_01948_));
 TAPCELL_X1 PHY_78 ();
 AOI22_X1 _06186_ (.A1(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[17][1] ),
    .A2(net79),
    .B1(net213),
    .B2(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[30][1] ),
    .ZN(_01950_));
 AOI22_X2 _06187_ (.A1(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[5][1] ),
    .A2(net134),
    .B1(net222),
    .B2(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[22][1] ),
    .ZN(_01951_));
 NAND4_X2 _06188_ (.A1(_01947_),
    .A2(_01948_),
    .A3(_01950_),
    .A4(_01951_),
    .ZN(_01952_));
 NOR4_X2 _06189_ (.A1(_01932_),
    .A2(_01938_),
    .A3(_01945_),
    .A4(_01952_),
    .ZN(_01953_));
 OAI21_X1 _06190_ (.A(_01295_),
    .B1(net130),
    .B2(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[0][1] ),
    .ZN(_01954_));
 OAI22_X2 _06191_ (.A1(_01925_),
    .A2(_01926_),
    .B1(_01953_),
    .B2(_01954_),
    .ZN(_01955_));
 AOI22_X1 _06192_ (.A1(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[23][1] ),
    .A2(net105),
    .B1(net197),
    .B2(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[19][1] ),
    .ZN(_01956_));
 AOI22_X1 _06193_ (.A1(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[8][1] ),
    .A2(net184),
    .B1(net206),
    .B2(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[13][1] ),
    .ZN(_01957_));
 TAPCELL_X1 PHY_77 ();
 AOI22_X1 _06195_ (.A1(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[17][1] ),
    .A2(net80),
    .B1(net264),
    .B2(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[18][1] ),
    .ZN(_01959_));
 AOI22_X2 _06196_ (.A1(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[12][1] ),
    .A2(net270),
    .B1(net243),
    .B2(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[2][1] ),
    .ZN(_01960_));
 NAND4_X2 _06197_ (.A1(_01956_),
    .A2(_01957_),
    .A3(_01959_),
    .A4(_01960_),
    .ZN(_01961_));
 AOI22_X1 _06198_ (.A1(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[5][1] ),
    .A2(net138),
    .B1(net85),
    .B2(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[14][1] ),
    .ZN(_01962_));
 AOI22_X1 _06199_ (.A1(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[3][1] ),
    .A2(net65),
    .B1(net247),
    .B2(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[20][1] ),
    .ZN(_01963_));
 AOI22_X1 _06200_ (.A1(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[9][1] ),
    .A2(net220),
    .B1(net210),
    .B2(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[30][1] ),
    .ZN(_01964_));
 NOR2_X1 _06201_ (.A1(net8),
    .A2(net9),
    .ZN(_01965_));
 TAPCELL_X1 PHY_76 ();
 NAND2_X1 _06203_ (.A1(net1),
    .A2(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[25][1] ),
    .ZN(_01967_));
 OAI22_X2 _06204_ (.A1(net1),
    .A2(_00985_),
    .B1(_01967_),
    .B2(_00992_),
    .ZN(_01968_));
 AOI22_X1 _06205_ (.A1(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[22][1] ),
    .A2(net225),
    .B1(_01965_),
    .B2(_01968_),
    .ZN(_01969_));
 NAND4_X1 _06206_ (.A1(_01962_),
    .A2(_01963_),
    .A3(_01964_),
    .A4(_01969_),
    .ZN(_01970_));
 AOI22_X1 _06207_ (.A1(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[28][1] ),
    .A2(net75),
    .B1(net82),
    .B2(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[21][1] ),
    .ZN(_01971_));
 AOI22_X1 _06208_ (.A1(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[27][1] ),
    .A2(net189),
    .B1(net96),
    .B2(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[31][1] ),
    .ZN(_01972_));
 AOI22_X1 _06209_ (.A1(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[26][1] ),
    .A2(net169),
    .B1(net143),
    .B2(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[29][1] ),
    .ZN(_01973_));
 AOI22_X1 _06210_ (.A1(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[16][1] ),
    .A2(net118),
    .B1(net259),
    .B2(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[1][1] ),
    .ZN(_01974_));
 NAND4_X1 _06211_ (.A1(_01971_),
    .A2(_01972_),
    .A3(_01973_),
    .A4(_01974_),
    .ZN(_01975_));
 AOI222_X2 _06212_ (.A1(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[15][1] ),
    .A2(net106),
    .B1(net164),
    .B2(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[6][1] ),
    .C1(net235),
    .C2(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[11][1] ),
    .ZN(_01976_));
 AOI22_X1 _06213_ (.A1(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[7][1] ),
    .A2(net67),
    .B1(net91),
    .B2(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[10][1] ),
    .ZN(_01977_));
 AOI22_X1 _06214_ (.A1(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[24][1] ),
    .A2(net72),
    .B1(net125),
    .B2(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[4][1] ),
    .ZN(_01978_));
 NAND3_X1 _06215_ (.A1(_01976_),
    .A2(_01977_),
    .A3(_01978_),
    .ZN(_01979_));
 NOR4_X2 _06216_ (.A1(_01961_),
    .A2(_01970_),
    .A3(_01975_),
    .A4(_01979_),
    .ZN(_01980_));
 OAI21_X1 _06217_ (.A(_01350_),
    .B1(_01064_),
    .B2(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[0][1] ),
    .ZN(_01981_));
 AOI22_X1 _06218_ (.A1(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[3][1] ),
    .A2(net65),
    .B1(net109),
    .B2(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[15][1] ),
    .ZN(_01982_));
 TAPCELL_X1 PHY_75 ();
 AOI22_X1 _06220_ (.A1(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[8][1] ),
    .A2(net182),
    .B1(net84),
    .B2(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[21][1] ),
    .ZN(_01984_));
 AOI22_X1 _06221_ (.A1(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[23][1] ),
    .A2(net98),
    .B1(net206),
    .B2(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[13][1] ),
    .ZN(_01985_));
 TAPCELL_X1 PHY_74 ();
 AOI22_X2 _06223_ (.A1(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[27][1] ),
    .A2(net191),
    .B1(net207),
    .B2(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[30][1] ),
    .ZN(_01987_));
 NAND4_X2 _06224_ (.A1(_01982_),
    .A2(_01984_),
    .A3(_01985_),
    .A4(_01987_),
    .ZN(_01988_));
 AOI22_X1 _06225_ (.A1(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[12][1] ),
    .A2(net266),
    .B1(net232),
    .B2(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[11][1] ),
    .ZN(_01989_));
 AOI22_X1 _06226_ (.A1(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[2][1] ),
    .A2(net243),
    .B1(net220),
    .B2(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[9][1] ),
    .ZN(_01990_));
 AOI22_X1 _06227_ (.A1(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[14][1] ),
    .A2(net86),
    .B1(net248),
    .B2(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[20][1] ),
    .ZN(_01991_));
 TAPCELL_X1 PHY_73 ();
 AOI21_X1 _06229_ (.A(_01119_),
    .B1(net264),
    .B2(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[18][1] ),
    .ZN(_01993_));
 NAND4_X1 _06230_ (.A1(_01989_),
    .A2(_01990_),
    .A3(_01991_),
    .A4(_01993_),
    .ZN(_01994_));
 AOI22_X1 _06231_ (.A1(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[25][1] ),
    .A2(net149),
    .B1(net140),
    .B2(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[29][1] ),
    .ZN(_01995_));
 AOI22_X1 _06232_ (.A1(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[31][1] ),
    .A2(_01149_),
    .B1(net223),
    .B2(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[22][1] ),
    .ZN(_01996_));
 AOI22_X1 _06233_ (.A1(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[16][1] ),
    .A2(net119),
    .B1(net128),
    .B2(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[4][1] ),
    .ZN(_01997_));
 TAPCELL_X1 PHY_72 ();
 AOI22_X2 _06235_ (.A1(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[7][1] ),
    .A2(net67),
    .B1(net91),
    .B2(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[10][1] ),
    .ZN(_01999_));
 NAND4_X2 _06236_ (.A1(_01995_),
    .A2(_01996_),
    .A3(_01997_),
    .A4(_01999_),
    .ZN(_02000_));
 AOI22_X1 _06237_ (.A1(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[17][1] ),
    .A2(net78),
    .B1(net72),
    .B2(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[24][1] ),
    .ZN(_02001_));
 AOI22_X1 _06238_ (.A1(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[1][1] ),
    .A2(net258),
    .B1(net197),
    .B2(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[19][1] ),
    .ZN(_02002_));
 AOI22_X1 _06239_ (.A1(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[28][1] ),
    .A2(net75),
    .B1(net164),
    .B2(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[6][1] ),
    .ZN(_02003_));
 AOI22_X1 _06240_ (.A1(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[26][1] ),
    .A2(net168),
    .B1(net136),
    .B2(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[5][1] ),
    .ZN(_02004_));
 NAND4_X2 _06241_ (.A1(_02001_),
    .A2(_02002_),
    .A3(_02003_),
    .A4(_02004_),
    .ZN(_02005_));
 NOR4_X2 _06242_ (.A1(_01988_),
    .A2(_01994_),
    .A3(_02000_),
    .A4(_02005_),
    .ZN(_02006_));
 OAI21_X1 _06243_ (.A(_00923_),
    .B1(_01064_),
    .B2(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[0][1] ),
    .ZN(_02007_));
 OAI22_X2 _06244_ (.A1(_01980_),
    .A2(_01981_),
    .B1(_02006_),
    .B2(_02007_),
    .ZN(_02008_));
 NOR4_X1 _06245_ (.A1(_01877_),
    .A2(_01902_),
    .A3(_01955_),
    .A4(_02008_),
    .ZN(_02009_));
 OAI21_X1 _06246_ (.A(_01731_),
    .B1(_01064_),
    .B2(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[0][1] ),
    .ZN(_02010_));
 INV_X1 _06247_ (.A(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[13][1] ),
    .ZN(_02011_));
 INV_X1 _06248_ (.A(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[24][1] ),
    .ZN(_02012_));
 OAI33_X1 _06249_ (.A1(_02011_),
    .A2(_01005_),
    .A3(_00948_),
    .B1(_00954_),
    .B2(_00979_),
    .B3(_02012_),
    .ZN(_02013_));
 AOI221_X1 _06250_ (.A(_02013_),
    .B1(_00975_),
    .B2(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[1][1] ),
    .C1(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[14][1] ),
    .C2(_00971_),
    .ZN(_02014_));
 INV_X1 _06251_ (.A(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[25][1] ),
    .ZN(_02015_));
 INV_X1 _06252_ (.A(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[22][1] ),
    .ZN(_02016_));
 OAI22_X1 _06253_ (.A1(_02015_),
    .A2(_01470_),
    .B1(_01216_),
    .B2(_02016_),
    .ZN(_02017_));
 AOI221_X1 _06254_ (.A(_02017_),
    .B1(net70),
    .B2(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[7][1] ),
    .C1(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[20][1] ),
    .C2(net244),
    .ZN(_02018_));
 INV_X1 _06255_ (.A(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[16][1] ),
    .ZN(_02019_));
 INV_X1 _06256_ (.A(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[26][1] ),
    .ZN(_02020_));
 OAI22_X1 _06257_ (.A1(_02019_),
    .A2(_01027_),
    .B1(_01203_),
    .B2(_02020_),
    .ZN(_02021_));
 AOI221_X1 _06258_ (.A(_02021_),
    .B1(net201),
    .B2(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[19][1] ),
    .C1(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[21][1] ),
    .C2(_00981_),
    .ZN(_02022_));
 INV_X1 _06259_ (.A(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[15][1] ),
    .ZN(_02023_));
 NAND2_X4 _06260_ (.A1(_00926_),
    .A2(_01026_),
    .ZN(_02024_));
 INV_X1 _06261_ (.A(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[18][1] ),
    .ZN(_02025_));
 OAI22_X1 _06262_ (.A1(_02023_),
    .A2(_01029_),
    .B1(_02024_),
    .B2(_02025_),
    .ZN(_02026_));
 AOI221_X1 _06263_ (.A(_02026_),
    .B1(_00989_),
    .B2(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[2][1] ),
    .C1(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[17][1] ),
    .C2(net81),
    .ZN(_02027_));
 AND4_X1 _06264_ (.A1(_02014_),
    .A2(_02018_),
    .A3(_02022_),
    .A4(_02027_),
    .ZN(_02028_));
 AOI22_X1 _06265_ (.A1(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[29][1] ),
    .A2(net146),
    .B1(net89),
    .B2(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[10][1] ),
    .ZN(_02029_));
 AOI22_X1 _06266_ (.A1(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[28][1] ),
    .A2(_01032_),
    .B1(net272),
    .B2(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[12][1] ),
    .ZN(_02030_));
 AOI22_X1 _06267_ (.A1(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[8][1] ),
    .A2(net183),
    .B1(net128),
    .B2(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[4][1] ),
    .ZN(_02031_));
 AOI22_X1 _06268_ (.A1(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[23][1] ),
    .A2(net99),
    .B1(net156),
    .B2(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[6][1] ),
    .ZN(_02032_));
 AND2_X1 _06269_ (.A1(_02031_),
    .A2(_02032_),
    .ZN(_02033_));
 AOI22_X1 _06270_ (.A1(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[27][1] ),
    .A2(_01021_),
    .B1(net211),
    .B2(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[30][1] ),
    .ZN(_02034_));
 NOR3_X4 _06271_ (.A1(_00953_),
    .A2(net10),
    .A3(net9),
    .ZN(_02035_));
 NOR2_X4 _06272_ (.A1(net1),
    .A2(_00978_),
    .ZN(_02036_));
 NAND3_X1 _06273_ (.A1(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[3][1] ),
    .A2(_02035_),
    .A3(_02036_),
    .ZN(_02037_));
 NAND2_X1 _06274_ (.A1(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[5][1] ),
    .A2(net139),
    .ZN(_02038_));
 INV_X1 _06275_ (.A(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[31][1] ),
    .ZN(_02039_));
 OAI33_X1 _06276_ (.A1(_02039_),
    .A2(_00960_),
    .A3(_01005_),
    .B1(_00948_),
    .B2(_00985_),
    .B3(net9),
    .ZN(_02040_));
 AOI221_X1 _06277_ (.A(_02040_),
    .B1(_00999_),
    .B2(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[9][1] ),
    .C1(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[11][1] ),
    .C2(net237),
    .ZN(_02041_));
 AND4_X1 _06278_ (.A1(_02034_),
    .A2(_02037_),
    .A3(_02038_),
    .A4(_02041_),
    .ZN(_02042_));
 AND4_X1 _06279_ (.A1(_02029_),
    .A2(_02030_),
    .A3(_02033_),
    .A4(_02042_),
    .ZN(_02043_));
 AOI21_X2 _06280_ (.A(_02010_),
    .B1(_02028_),
    .B2(_02043_),
    .ZN(_02044_));
 NOR2_X1 _06281_ (.A1(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[0][1] ),
    .A2(net130),
    .ZN(_02045_));
 NOR4_X1 _06282_ (.A1(net4),
    .A2(net5),
    .A3(_01349_),
    .A4(_02045_),
    .ZN(_02046_));
 AOI22_X1 _06283_ (.A1(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[2][1] ),
    .A2(net239),
    .B1(net221),
    .B2(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[9][1] ),
    .ZN(_02047_));
 AOI22_X1 _06284_ (.A1(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[18][1] ),
    .A2(_00964_),
    .B1(net200),
    .B2(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[19][1] ),
    .ZN(_02048_));
 AOI22_X1 _06285_ (.A1(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[8][1] ),
    .A2(net177),
    .B1(net89),
    .B2(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[10][1] ),
    .ZN(_02049_));
 AOI22_X1 _06286_ (.A1(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[17][1] ),
    .A2(net81),
    .B1(net186),
    .B2(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[27][1] ),
    .ZN(_02050_));
 NAND4_X1 _06287_ (.A1(_02047_),
    .A2(_02048_),
    .A3(_02049_),
    .A4(_02050_),
    .ZN(_02051_));
 AOI22_X1 _06288_ (.A1(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[6][1] ),
    .A2(net159),
    .B1(net216),
    .B2(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[30][1] ),
    .ZN(_02052_));
 AOI22_X1 _06289_ (.A1(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[26][1] ),
    .A2(net167),
    .B1(net274),
    .B2(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[12][1] ),
    .ZN(_02053_));
 MUX2_X1 _06290_ (.A(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[5][1] ),
    .B(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[21][1] ),
    .S(net1),
    .Z(_02054_));
 AOI221_X1 _06291_ (.A(net115),
    .B1(_01597_),
    .B2(_02054_),
    .C1(net151),
    .C2(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[25][1] ),
    .ZN(_02055_));
 NAND3_X1 _06292_ (.A1(_02052_),
    .A2(_02053_),
    .A3(_02055_),
    .ZN(_02056_));
 AOI22_X1 _06293_ (.A1(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[23][1] ),
    .A2(_01144_),
    .B1(_01032_),
    .B2(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[28][1] ),
    .ZN(_02057_));
 AOI22_X1 _06294_ (.A1(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[16][1] ),
    .A2(net121),
    .B1(net262),
    .B2(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[1][1] ),
    .ZN(_02058_));
 AOI22_X1 _06295_ (.A1(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[7][1] ),
    .A2(net70),
    .B1(net88),
    .B2(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[14][1] ),
    .ZN(_02059_));
 AOI22_X1 _06296_ (.A1(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[31][1] ),
    .A2(net94),
    .B1(net244),
    .B2(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[20][1] ),
    .ZN(_02060_));
 NAND4_X1 _06297_ (.A1(_02057_),
    .A2(_02058_),
    .A3(_02059_),
    .A4(_02060_),
    .ZN(_02061_));
 AOI22_X1 _06298_ (.A1(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[29][1] ),
    .A2(net141),
    .B1(_01007_),
    .B2(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[13][1] ),
    .ZN(_02062_));
 AOI22_X1 _06299_ (.A1(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[4][1] ),
    .A2(net129),
    .B1(_00993_),
    .B2(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[11][1] ),
    .ZN(_02063_));
 AOI22_X1 _06300_ (.A1(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[3][1] ),
    .A2(net63),
    .B1(_00996_),
    .B2(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[22][1] ),
    .ZN(_02064_));
 AOI22_X1 _06301_ (.A1(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[15][1] ),
    .A2(net111),
    .B1(_01059_),
    .B2(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[24][1] ),
    .ZN(_02065_));
 NAND4_X1 _06302_ (.A1(_02062_),
    .A2(_02063_),
    .A3(_02064_),
    .A4(_02065_),
    .ZN(_02066_));
 OR4_X2 _06303_ (.A1(_02051_),
    .A2(_02056_),
    .A3(_02061_),
    .A4(_02066_),
    .ZN(_02067_));
 AOI21_X1 _06304_ (.A(_02044_),
    .B1(_02046_),
    .B2(_02067_),
    .ZN(_02068_));
 AOI22_X1 _06305_ (.A1(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[17][1] ),
    .A2(net79),
    .B1(net66),
    .B2(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[3][1] ),
    .ZN(_02069_));
 AOI22_X1 _06306_ (.A1(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[6][1] ),
    .A2(net162),
    .B1(net222),
    .B2(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[22][1] ),
    .ZN(_02070_));
 TAPCELL_X1 PHY_71 ();
 AOI22_X1 _06308_ (.A1(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[31][1] ),
    .A2(net93),
    .B1(net193),
    .B2(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[19][1] ),
    .ZN(_02072_));
 AOI22_X1 _06309_ (.A1(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[16][1] ),
    .A2(net116),
    .B1(net263),
    .B2(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[18][1] ),
    .ZN(_02073_));
 NAND4_X1 _06310_ (.A1(_02069_),
    .A2(_02070_),
    .A3(_02072_),
    .A4(_02073_),
    .ZN(_02074_));
 AOI22_X1 _06311_ (.A1(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[23][1] ),
    .A2(net104),
    .B1(net250),
    .B2(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[20][1] ),
    .ZN(_02075_));
 AOI22_X1 _06312_ (.A1(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[15][1] ),
    .A2(net108),
    .B1(net123),
    .B2(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[4][1] ),
    .ZN(_02076_));
 MUX2_X1 _06313_ (.A(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[12][1] ),
    .B(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[14][1] ),
    .S(net8),
    .Z(_02077_));
 AOI221_X1 _06314_ (.A(net114),
    .B1(net92),
    .B2(_02077_),
    .C1(net240),
    .C2(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[2][1] ),
    .ZN(_02078_));
 NAND3_X1 _06315_ (.A1(_02075_),
    .A2(_02076_),
    .A3(_02078_),
    .ZN(_02079_));
 AOI22_X1 _06316_ (.A1(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[24][1] ),
    .A2(net71),
    .B1(net255),
    .B2(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[1][1] ),
    .ZN(_02080_));
 AOI22_X1 _06317_ (.A1(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[25][1] ),
    .A2(net152),
    .B1(net217),
    .B2(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[9][1] ),
    .ZN(_02081_));
 AOI22_X1 _06318_ (.A1(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[27][1] ),
    .A2(net188),
    .B1(net204),
    .B2(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[13][1] ),
    .ZN(_02082_));
 AOI22_X1 _06319_ (.A1(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[26][1] ),
    .A2(net173),
    .B1(net83),
    .B2(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[21][1] ),
    .ZN(_02083_));
 NAND4_X1 _06320_ (.A1(_02080_),
    .A2(_02081_),
    .A3(_02082_),
    .A4(_02083_),
    .ZN(_02084_));
 AOI22_X1 _06321_ (.A1(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[28][1] ),
    .A2(net76),
    .B1(net180),
    .B2(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[8][1] ),
    .ZN(_02085_));
 AOI22_X1 _06322_ (.A1(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[5][1] ),
    .A2(net131),
    .B1(net68),
    .B2(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[7][1] ),
    .ZN(_02086_));
 AOI22_X1 _06323_ (.A1(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[29][1] ),
    .A2(net144),
    .B1(net233),
    .B2(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[11][1] ),
    .ZN(_02087_));
 AOI22_X1 _06324_ (.A1(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[10][1] ),
    .A2(net90),
    .B1(net208),
    .B2(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[30][1] ),
    .ZN(_02088_));
 NAND4_X1 _06325_ (.A1(_02085_),
    .A2(_02086_),
    .A3(_02087_),
    .A4(_02088_),
    .ZN(_02089_));
 OR4_X1 _06326_ (.A1(_02074_),
    .A2(_02079_),
    .A3(_02084_),
    .A4(_02089_),
    .ZN(_02090_));
 NOR2_X1 _06327_ (.A1(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[0][1] ),
    .A2(net130),
    .ZN(_02091_));
 NOR3_X1 _06328_ (.A1(_00922_),
    .A2(_01349_),
    .A3(_02091_),
    .ZN(_02092_));
 AOI22_X1 _06329_ (.A1(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[17][1] ),
    .A2(net78),
    .B1(net212),
    .B2(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[30][1] ),
    .ZN(_02093_));
 AOI22_X1 _06330_ (.A1(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[15][1] ),
    .A2(net108),
    .B1(net260),
    .B2(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[1][1] ),
    .ZN(_02094_));
 AOI22_X1 _06331_ (.A1(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[28][1] ),
    .A2(net77),
    .B1(net271),
    .B2(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[12][1] ),
    .ZN(_02095_));
 AOI22_X1 _06332_ (.A1(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[8][1] ),
    .A2(_01034_),
    .B1(net72),
    .B2(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[24][1] ),
    .ZN(_02096_));
 NAND4_X1 _06333_ (.A1(_02093_),
    .A2(_02094_),
    .A3(_02095_),
    .A4(_02096_),
    .ZN(_02097_));
 AOI22_X1 _06334_ (.A1(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[3][1] ),
    .A2(net65),
    .B1(net235),
    .B2(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[11][1] ),
    .ZN(_02098_));
 AOI22_X1 _06335_ (.A1(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[16][1] ),
    .A2(net118),
    .B1(net86),
    .B2(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[14][1] ),
    .ZN(_02099_));
 AOI22_X1 _06336_ (.A1(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[29][1] ),
    .A2(net143),
    .B1(net249),
    .B2(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[20][1] ),
    .ZN(_02100_));
 AOI21_X1 _06337_ (.A(net114),
    .B1(net105),
    .B2(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[23][1] ),
    .ZN(_02101_));
 NAND4_X1 _06338_ (.A1(_02098_),
    .A2(_02099_),
    .A3(_02100_),
    .A4(_02101_),
    .ZN(_02102_));
 AOI22_X1 _06339_ (.A1(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[26][1] ),
    .A2(_01038_),
    .B1(net220),
    .B2(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[9][1] ),
    .ZN(_02103_));
 AOI22_X1 _06340_ (.A1(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[27][1] ),
    .A2(net191),
    .B1(net96),
    .B2(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[31][1] ),
    .ZN(_02104_));
 AOI22_X1 _06341_ (.A1(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[5][1] ),
    .A2(net138),
    .B1(net84),
    .B2(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[21][1] ),
    .ZN(_02105_));
 AOI22_X1 _06342_ (.A1(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[25][1] ),
    .A2(net155),
    .B1(net241),
    .B2(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[2][1] ),
    .ZN(_02106_));
 NAND4_X1 _06343_ (.A1(_02103_),
    .A2(_02104_),
    .A3(_02105_),
    .A4(_02106_),
    .ZN(_02107_));
 AOI22_X1 _06344_ (.A1(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[7][1] ),
    .A2(net68),
    .B1(net265),
    .B2(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[18][1] ),
    .ZN(_02108_));
 AOI22_X1 _06345_ (.A1(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[6][1] ),
    .A2(net164),
    .B1(net91),
    .B2(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[10][1] ),
    .ZN(_02109_));
 AOI22_X1 _06346_ (.A1(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[4][1] ),
    .A2(net125),
    .B1(net224),
    .B2(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[22][1] ),
    .ZN(_02110_));
 AOI22_X1 _06347_ (.A1(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[13][1] ),
    .A2(net205),
    .B1(net196),
    .B2(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[19][1] ),
    .ZN(_02111_));
 NAND4_X1 _06348_ (.A1(_02108_),
    .A2(_02109_),
    .A3(_02110_),
    .A4(_02111_),
    .ZN(_02112_));
 OR4_X1 _06349_ (.A1(_02097_),
    .A2(_02102_),
    .A3(_02107_),
    .A4(_02112_),
    .ZN(_02113_));
 NOR2_X1 _06350_ (.A1(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[0][1] ),
    .A2(net130),
    .ZN(_02114_));
 NOR3_X1 _06351_ (.A1(_01163_),
    .A2(_01407_),
    .A3(_02114_),
    .ZN(_02115_));
 AOI22_X1 _06352_ (.A1(_02090_),
    .A2(_02092_),
    .B1(_02113_),
    .B2(_02115_),
    .ZN(_02116_));
 AOI22_X1 _06353_ (.A1(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[5][1] ),
    .A2(net134),
    .B1(net242),
    .B2(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[2][1] ),
    .ZN(_02117_));
 AOI22_X1 _06354_ (.A1(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[31][1] ),
    .A2(net93),
    .B1(net226),
    .B2(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[22][1] ),
    .ZN(_02118_));
 AOI22_X1 _06355_ (.A1(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[14][1] ),
    .A2(net87),
    .B1(net212),
    .B2(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[30][1] ),
    .ZN(_02119_));
 AOI22_X1 _06356_ (.A1(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[6][1] ),
    .A2(net163),
    .B1(net269),
    .B2(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[12][1] ),
    .ZN(_02120_));
 NAND4_X1 _06357_ (.A1(_02117_),
    .A2(_02118_),
    .A3(_02119_),
    .A4(_02120_),
    .ZN(_02121_));
 AOI22_X1 _06358_ (.A1(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[16][1] ),
    .A2(net117),
    .B1(net77),
    .B2(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[28][1] ),
    .ZN(_02122_));
 AOI22_X1 _06359_ (.A1(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[23][1] ),
    .A2(net101),
    .B1(net90),
    .B2(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[10][1] ),
    .ZN(_02123_));
 AOI22_X1 _06360_ (.A1(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[29][1] ),
    .A2(net144),
    .B1(net260),
    .B2(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[1][1] ),
    .ZN(_02124_));
 AOI21_X1 _06361_ (.A(net114),
    .B1(net263),
    .B2(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[18][1] ),
    .ZN(_02125_));
 NAND4_X1 _06362_ (.A1(_02122_),
    .A2(_02123_),
    .A3(_02124_),
    .A4(_02125_),
    .ZN(_02126_));
 AOI22_X1 _06363_ (.A1(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[15][1] ),
    .A2(net108),
    .B1(net203),
    .B2(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[13][1] ),
    .ZN(_02127_));
 AOI22_X1 _06364_ (.A1(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[26][1] ),
    .A2(net175),
    .B1(net245),
    .B2(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[20][1] ),
    .ZN(_02128_));
 AOI22_X1 _06365_ (.A1(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[27][1] ),
    .A2(net188),
    .B1(net218),
    .B2(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[9][1] ),
    .ZN(_02129_));
 AOI22_X1 _06366_ (.A1(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[25][1] ),
    .A2(net148),
    .B1(net83),
    .B2(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[21][1] ),
    .ZN(_02130_));
 NAND4_X1 _06367_ (.A1(_02127_),
    .A2(_02128_),
    .A3(_02129_),
    .A4(_02130_),
    .ZN(_02131_));
 AOI22_X1 _06368_ (.A1(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[17][1] ),
    .A2(net79),
    .B1(net236),
    .B2(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[11][1] ),
    .ZN(_02132_));
 AOI22_X1 _06369_ (.A1(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[8][1] ),
    .A2(net180),
    .B1(net126),
    .B2(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[4][1] ),
    .ZN(_02133_));
 AOI22_X1 _06370_ (.A1(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[24][1] ),
    .A2(net71),
    .B1(net193),
    .B2(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[19][1] ),
    .ZN(_02134_));
 AOI22_X1 _06371_ (.A1(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[3][1] ),
    .A2(net66),
    .B1(net68),
    .B2(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[7][1] ),
    .ZN(_02135_));
 NAND4_X1 _06372_ (.A1(_02132_),
    .A2(_02133_),
    .A3(_02134_),
    .A4(_02135_),
    .ZN(_02136_));
 OR4_X1 _06373_ (.A1(_02121_),
    .A2(_02126_),
    .A3(_02131_),
    .A4(_02136_),
    .ZN(_02137_));
 OAI21_X1 _06374_ (.A(_01700_),
    .B1(net130),
    .B2(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[0][1] ),
    .ZN(_02138_));
 INV_X1 _06375_ (.A(_02138_),
    .ZN(_02139_));
 AOI22_X1 _06376_ (.A1(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[7][1] ),
    .A2(net70),
    .B1(net129),
    .B2(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[4][1] ),
    .ZN(_02140_));
 AOI22_X1 _06377_ (.A1(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[21][1] ),
    .A2(_00981_),
    .B1(net215),
    .B2(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[30][1] ),
    .ZN(_02141_));
 AOI22_X1 _06378_ (.A1(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[27][1] ),
    .A2(net186),
    .B1(_01149_),
    .B2(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[31][1] ),
    .ZN(_02142_));
 AOI22_X1 _06379_ (.A1(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[3][1] ),
    .A2(net63),
    .B1(net156),
    .B2(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[6][1] ),
    .ZN(_02143_));
 NAND4_X1 _06380_ (.A1(_02140_),
    .A2(_02141_),
    .A3(_02142_),
    .A4(_02143_),
    .ZN(_02144_));
 AOI222_X2 _06381_ (.A1(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[15][1] ),
    .A2(net111),
    .B1(net135),
    .B2(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[5][1] ),
    .C1(net244),
    .C2(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[20][1] ),
    .ZN(_02145_));
 AOI22_X1 _06382_ (.A1(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[28][1] ),
    .A2(_01032_),
    .B1(_00964_),
    .B2(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[18][1] ),
    .ZN(_02146_));
 AOI22_X1 _06383_ (.A1(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[22][1] ),
    .A2(_00996_),
    .B1(_01007_),
    .B2(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[13][1] ),
    .ZN(_02147_));
 NAND3_X1 _06384_ (.A1(_02145_),
    .A2(_02146_),
    .A3(_02147_),
    .ZN(_02148_));
 AOI221_X1 _06385_ (.A(net115),
    .B1(_00975_),
    .B2(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[1][1] ),
    .C1(_00989_),
    .C2(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[2][1] ),
    .ZN(_02149_));
 AOI22_X1 _06386_ (.A1(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[17][1] ),
    .A2(net81),
    .B1(net151),
    .B2(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[25][1] ),
    .ZN(_02150_));
 AOI22_X1 _06387_ (.A1(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[16][1] ),
    .A2(net121),
    .B1(net88),
    .B2(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[14][1] ),
    .ZN(_02151_));
 AOI22_X1 _06388_ (.A1(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[23][1] ),
    .A2(_01144_),
    .B1(net176),
    .B2(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[8][1] ),
    .ZN(_02152_));
 NAND4_X1 _06389_ (.A1(_02149_),
    .A2(_02150_),
    .A3(_02151_),
    .A4(_02152_),
    .ZN(_02153_));
 AOI22_X1 _06390_ (.A1(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[12][1] ),
    .A2(net274),
    .B1(net89),
    .B2(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[10][1] ),
    .ZN(_02154_));
 AOI22_X1 _06391_ (.A1(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[26][1] ),
    .A2(net167),
    .B1(_01050_),
    .B2(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[29][1] ),
    .ZN(_02155_));
 AOI22_X1 _06392_ (.A1(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[24][1] ),
    .A2(_01059_),
    .B1(net221),
    .B2(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[9][1] ),
    .ZN(_02156_));
 AOI22_X1 _06393_ (.A1(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[11][1] ),
    .A2(net231),
    .B1(net200),
    .B2(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[19][1] ),
    .ZN(_02157_));
 NAND4_X1 _06394_ (.A1(_02154_),
    .A2(_02155_),
    .A3(_02156_),
    .A4(_02157_),
    .ZN(_02158_));
 OR4_X2 _06395_ (.A1(_02144_),
    .A2(_02148_),
    .A3(_02153_),
    .A4(_02158_),
    .ZN(_02159_));
 OAI21_X1 _06396_ (.A(_01502_),
    .B1(net130),
    .B2(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[0][1] ),
    .ZN(_02160_));
 INV_X1 _06397_ (.A(_02160_),
    .ZN(_02161_));
 AOI22_X1 _06398_ (.A1(_02137_),
    .A2(_02139_),
    .B1(_02159_),
    .B2(_02161_),
    .ZN(_02162_));
 AOI22_X1 _06399_ (.A1(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[17][1] ),
    .A2(net78),
    .B1(net86),
    .B2(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[14][1] ),
    .ZN(_02163_));
 AOI22_X1 _06400_ (.A1(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[29][1] ),
    .A2(net140),
    .B1(net248),
    .B2(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[20][1] ),
    .ZN(_02164_));
 AOI22_X1 _06401_ (.A1(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[27][1] ),
    .A2(net189),
    .B1(net149),
    .B2(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[25][1] ),
    .ZN(_02165_));
 AOI22_X1 _06402_ (.A1(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[26][1] ),
    .A2(net168),
    .B1(net136),
    .B2(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[5][1] ),
    .ZN(_02166_));
 NAND4_X1 _06403_ (.A1(_02163_),
    .A2(_02164_),
    .A3(_02165_),
    .A4(_02166_),
    .ZN(_02167_));
 AOI22_X1 _06404_ (.A1(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[16][1] ),
    .A2(net118),
    .B1(net82),
    .B2(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[21][1] ),
    .ZN(_02168_));
 AOI22_X1 _06405_ (.A1(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[6][1] ),
    .A2(net161),
    .B1(net257),
    .B2(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[1][1] ),
    .ZN(_02169_));
 AOI22_X1 _06406_ (.A1(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[15][1] ),
    .A2(net106),
    .B1(net75),
    .B2(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[28][1] ),
    .ZN(_02170_));
 AOI21_X1 _06407_ (.A(net113),
    .B1(net220),
    .B2(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[9][1] ),
    .ZN(_02171_));
 NAND4_X2 _06408_ (.A1(_02168_),
    .A2(_02169_),
    .A3(_02170_),
    .A4(_02171_),
    .ZN(_02172_));
 AOI22_X1 _06409_ (.A1(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[18][1] ),
    .A2(net264),
    .B1(net197),
    .B2(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[19][1] ),
    .ZN(_02173_));
 AOI22_X1 _06410_ (.A1(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[23][1] ),
    .A2(net98),
    .B1(net232),
    .B2(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[11][1] ),
    .ZN(_02174_));
 AOI22_X1 _06411_ (.A1(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[2][1] ),
    .A2(net243),
    .B1(net223),
    .B2(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[22][1] ),
    .ZN(_02175_));
 AOI22_X1 _06412_ (.A1(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[8][1] ),
    .A2(net183),
    .B1(net206),
    .B2(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[13][1] ),
    .ZN(_02176_));
 NAND4_X1 _06413_ (.A1(_02173_),
    .A2(_02174_),
    .A3(_02175_),
    .A4(_02176_),
    .ZN(_02177_));
 AOI22_X1 _06414_ (.A1(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[4][1] ),
    .A2(net125),
    .B1(net210),
    .B2(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[30][1] ),
    .ZN(_02178_));
 AOI22_X1 _06415_ (.A1(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[31][1] ),
    .A2(net96),
    .B1(net91),
    .B2(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[10][1] ),
    .ZN(_02179_));
 AOI22_X1 _06416_ (.A1(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[3][1] ),
    .A2(net65),
    .B1(net266),
    .B2(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[12][1] ),
    .ZN(_02180_));
 AOI22_X1 _06417_ (.A1(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[24][1] ),
    .A2(net72),
    .B1(net67),
    .B2(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[7][1] ),
    .ZN(_02181_));
 NAND4_X1 _06418_ (.A1(_02178_),
    .A2(_02179_),
    .A3(_02180_),
    .A4(_02181_),
    .ZN(_02182_));
 OR4_X2 _06419_ (.A1(_02167_),
    .A2(_02172_),
    .A3(_02177_),
    .A4(_02182_),
    .ZN(_02183_));
 OAI21_X1 _06420_ (.A(_01164_),
    .B1(net130),
    .B2(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[0][1] ),
    .ZN(_02184_));
 INV_X1 _06421_ (.A(_02184_),
    .ZN(_02185_));
 AOI22_X1 _06422_ (.A1(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[26][1] ),
    .A2(net170),
    .B1(net96),
    .B2(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[31][1] ),
    .ZN(_02186_));
 AOI22_X1 _06423_ (.A1(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[29][1] ),
    .A2(net145),
    .B1(net82),
    .B2(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[21][1] ),
    .ZN(_02187_));
 AOI22_X1 _06424_ (.A1(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[12][1] ),
    .A2(net271),
    .B1(net209),
    .B2(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[30][1] ),
    .ZN(_02188_));
 AOI22_X1 _06425_ (.A1(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[14][1] ),
    .A2(net85),
    .B1(net234),
    .B2(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[11][1] ),
    .ZN(_02189_));
 NAND4_X1 _06426_ (.A1(_02186_),
    .A2(_02187_),
    .A3(_02188_),
    .A4(_02189_),
    .ZN(_02190_));
 AOI22_X1 _06427_ (.A1(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[8][1] ),
    .A2(net184),
    .B1(net259),
    .B2(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[1][1] ),
    .ZN(_02191_));
 AOI22_X1 _06428_ (.A1(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[25][1] ),
    .A2(net154),
    .B1(net124),
    .B2(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[4][1] ),
    .ZN(_02192_));
 AOI22_X1 _06429_ (.A1(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[5][1] ),
    .A2(net137),
    .B1(net241),
    .B2(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[2][1] ),
    .ZN(_02193_));
 AOI21_X1 _06430_ (.A(net113),
    .B1(net219),
    .B2(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[9][1] ),
    .ZN(_02194_));
 NAND4_X1 _06431_ (.A1(_02191_),
    .A2(_02192_),
    .A3(_02193_),
    .A4(_02194_),
    .ZN(_02195_));
 AOI22_X1 _06432_ (.A1(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[23][1] ),
    .A2(net101),
    .B1(net265),
    .B2(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[18][1] ),
    .ZN(_02196_));
 AOI22_X1 _06433_ (.A1(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[17][1] ),
    .A2(net80),
    .B1(net224),
    .B2(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[22][1] ),
    .ZN(_02197_));
 AOI22_X1 _06434_ (.A1(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[7][1] ),
    .A2(net67),
    .B1(net90),
    .B2(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[10][1] ),
    .ZN(_02198_));
 AOI22_X1 _06435_ (.A1(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[24][1] ),
    .A2(net74),
    .B1(net249),
    .B2(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[20][1] ),
    .ZN(_02199_));
 NAND4_X1 _06436_ (.A1(_02196_),
    .A2(_02197_),
    .A3(_02198_),
    .A4(_02199_),
    .ZN(_02200_));
 AOI22_X1 _06437_ (.A1(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[15][1] ),
    .A2(net106),
    .B1(net195),
    .B2(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[19][1] ),
    .ZN(_02201_));
 AOI22_X1 _06438_ (.A1(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[3][1] ),
    .A2(net64),
    .B1(net118),
    .B2(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[16][1] ),
    .ZN(_02202_));
 AOI22_X1 _06439_ (.A1(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[28][1] ),
    .A2(net75),
    .B1(net163),
    .B2(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[6][1] ),
    .ZN(_02203_));
 AOI22_X1 _06440_ (.A1(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[27][1] ),
    .A2(net189),
    .B1(net205),
    .B2(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[13][1] ),
    .ZN(_02204_));
 NAND4_X1 _06441_ (.A1(_02201_),
    .A2(_02202_),
    .A3(_02203_),
    .A4(_02204_),
    .ZN(_02205_));
 OR4_X1 _06442_ (.A1(_02190_),
    .A2(_02195_),
    .A3(_02200_),
    .A4(_02205_),
    .ZN(_02206_));
 OAI21_X1 _06443_ (.A(_01169_),
    .B1(net130),
    .B2(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[0][1] ),
    .ZN(_02207_));
 INV_X1 _06444_ (.A(_02207_),
    .ZN(_02208_));
 AOI22_X1 _06445_ (.A1(_02183_),
    .A2(_02185_),
    .B1(_02206_),
    .B2(_02208_),
    .ZN(_02209_));
 AND4_X1 _06446_ (.A1(_02068_),
    .A2(_02116_),
    .A3(_02162_),
    .A4(_02209_),
    .ZN(_02210_));
 AOI22_X1 _06447_ (.A1(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[26][1] ),
    .A2(net173),
    .B1(net90),
    .B2(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[10][1] ),
    .ZN(_02211_));
 AOI22_X1 _06448_ (.A1(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[3][1] ),
    .A2(net64),
    .B1(net85),
    .B2(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[14][1] ),
    .ZN(_02212_));
 AOI22_X1 _06449_ (.A1(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[8][1] ),
    .A2(net179),
    .B1(net250),
    .B2(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[20][1] ),
    .ZN(_02213_));
 AOI22_X1 _06450_ (.A1(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[27][1] ),
    .A2(net190),
    .B1(net153),
    .B2(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[25][1] ),
    .ZN(_02214_));
 NAND4_X1 _06451_ (.A1(_02211_),
    .A2(_02212_),
    .A3(_02213_),
    .A4(_02214_),
    .ZN(_02215_));
 AOI22_X1 _06452_ (.A1(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[23][1] ),
    .A2(net100),
    .B1(net116),
    .B2(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[16][1] ),
    .ZN(_02216_));
 AOI22_X1 _06453_ (.A1(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[17][1] ),
    .A2(net79),
    .B1(net217),
    .B2(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[9][1] ),
    .ZN(_02217_));
 AOI22_X1 _06454_ (.A1(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[30][1] ),
    .A2(net208),
    .B1(net204),
    .B2(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[13][1] ),
    .ZN(_02218_));
 AOI21_X1 _06455_ (.A(net113),
    .B1(net194),
    .B2(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[19][1] ),
    .ZN(_02219_));
 NAND4_X1 _06456_ (.A1(_02216_),
    .A2(_02217_),
    .A3(_02218_),
    .A4(_02219_),
    .ZN(_02220_));
 AOI22_X1 _06457_ (.A1(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[15][1] ),
    .A2(net107),
    .B1(net93),
    .B2(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[31][1] ),
    .ZN(_02221_));
 AOI22_X1 _06458_ (.A1(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[5][1] ),
    .A2(net131),
    .B1(net82),
    .B2(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[21][1] ),
    .ZN(_02222_));
 AOI22_X1 _06459_ (.A1(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[29][1] ),
    .A2(net142),
    .B1(net255),
    .B2(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[1][1] ),
    .ZN(_02223_));
 AOI22_X1 _06460_ (.A1(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[7][1] ),
    .A2(net68),
    .B1(net233),
    .B2(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[11][1] ),
    .ZN(_02224_));
 NAND4_X1 _06461_ (.A1(_02221_),
    .A2(_02222_),
    .A3(_02223_),
    .A4(_02224_),
    .ZN(_02225_));
 AOI22_X1 _06462_ (.A1(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[24][1] ),
    .A2(net71),
    .B1(net240),
    .B2(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[2][1] ),
    .ZN(_02226_));
 AOI22_X1 _06463_ (.A1(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[4][1] ),
    .A2(net123),
    .B1(net263),
    .B2(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[18][1] ),
    .ZN(_02227_));
 AOI22_X1 _06464_ (.A1(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[12][1] ),
    .A2(net267),
    .B1(net226),
    .B2(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[22][1] ),
    .ZN(_02228_));
 AOI22_X1 _06465_ (.A1(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[28][1] ),
    .A2(net77),
    .B1(net162),
    .B2(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[6][1] ),
    .ZN(_02229_));
 NAND4_X1 _06466_ (.A1(_02226_),
    .A2(_02227_),
    .A3(_02228_),
    .A4(_02229_),
    .ZN(_02230_));
 OR4_X2 _06467_ (.A1(_02215_),
    .A2(_02220_),
    .A3(_02225_),
    .A4(_02230_),
    .ZN(_02231_));
 OAI21_X1 _06468_ (.A(_02231_),
    .B1(net130),
    .B2(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[0][1] ),
    .ZN(_02232_));
 AOI221_X2 _06469_ (.A(_00907_),
    .B1(_02009_),
    .B2(_02210_),
    .C1(_02232_),
    .C2(_01820_),
    .ZN(\rdata_o_n[1] ));
 TAPCELL_X1 PHY_70 ();
 AOI22_X1 _06471_ (.A1(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[31][2] ),
    .A2(net96),
    .B1(net225),
    .B2(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[22][2] ),
    .ZN(_02234_));
 AOI22_X1 _06472_ (.A1(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[4][2] ),
    .A2(net125),
    .B1(net241),
    .B2(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[2][2] ),
    .ZN(_02235_));
 AND2_X1 _06473_ (.A1(_02234_),
    .A2(_02235_),
    .ZN(_02236_));
 INV_X1 _06474_ (.A(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[16][2] ),
    .ZN(_02237_));
 NAND4_X4 _06475_ (.A1(net7),
    .A2(_00944_),
    .A3(net9),
    .A4(_00939_),
    .ZN(_02238_));
 INV_X1 _06476_ (.A(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[5][2] ),
    .ZN(_02239_));
 OAI22_X1 _06477_ (.A1(_02237_),
    .A2(_01027_),
    .B1(_02238_),
    .B2(_02239_),
    .ZN(_02240_));
 AOI221_X1 _06478_ (.A(_02240_),
    .B1(net235),
    .B2(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[11][2] ),
    .C1(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[28][2] ),
    .C2(net75),
    .ZN(_02241_));
 INV_X1 _06479_ (.A(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[17][2] ),
    .ZN(_02242_));
 INV_X1 _06480_ (.A(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[30][2] ),
    .ZN(_02243_));
 OAI33_X1 _06481_ (.A1(_02242_),
    .A2(_01015_),
    .A3(_00979_),
    .B1(_00960_),
    .B2(_00970_),
    .B3(_02243_),
    .ZN(_02244_));
 AOI221_X1 _06482_ (.A(_02244_),
    .B1(net91),
    .B2(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[10][2] ),
    .C1(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[21][2] ),
    .C2(net82),
    .ZN(_02245_));
 INV_X1 _06483_ (.A(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[12][2] ),
    .ZN(_02246_));
 OAI21_X1 _06484_ (.A(_01064_),
    .B1(_01426_),
    .B2(_02246_),
    .ZN(_02247_));
 AOI221_X1 _06485_ (.A(_02247_),
    .B1(net67),
    .B2(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[7][2] ),
    .C1(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[24][2] ),
    .C2(net72),
    .ZN(_02248_));
 NAND4_X1 _06486_ (.A1(_02236_),
    .A2(_02241_),
    .A3(_02245_),
    .A4(_02248_),
    .ZN(_02249_));
 AOI22_X1 _06487_ (.A1(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[6][2] ),
    .A2(net161),
    .B1(net257),
    .B2(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[1][2] ),
    .ZN(_02250_));
 AOI22_X1 _06488_ (.A1(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[27][2] ),
    .A2(net189),
    .B1(net103),
    .B2(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[23][2] ),
    .ZN(_02251_));
 AOI22_X1 _06489_ (.A1(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[8][2] ),
    .A2(net184),
    .B1(net205),
    .B2(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[13][2] ),
    .ZN(_02252_));
 AOI22_X1 _06490_ (.A1(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[29][2] ),
    .A2(net143),
    .B1(net265),
    .B2(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[18][2] ),
    .ZN(_02253_));
 AND4_X1 _06491_ (.A1(_02250_),
    .A2(_02251_),
    .A3(_02252_),
    .A4(_02253_),
    .ZN(_02254_));
 AOI22_X1 _06492_ (.A1(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[14][2] ),
    .A2(net85),
    .B1(net247),
    .B2(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[20][2] ),
    .ZN(_02255_));
 AOI22_X1 _06493_ (.A1(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[3][2] ),
    .A2(net64),
    .B1(net220),
    .B2(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[9][2] ),
    .ZN(_02256_));
 AOI22_X1 _06494_ (.A1(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[26][2] ),
    .A2(net169),
    .B1(_01009_),
    .B2(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[19][2] ),
    .ZN(_02257_));
 TAPCELL_X1 PHY_69 ();
 AOI22_X1 _06496_ (.A1(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[15][2] ),
    .A2(net106),
    .B1(net154),
    .B2(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[25][2] ),
    .ZN(_02259_));
 AND2_X1 _06497_ (.A1(_02257_),
    .A2(_02259_),
    .ZN(_02260_));
 NAND4_X2 _06498_ (.A1(_02254_),
    .A2(_02255_),
    .A3(_02256_),
    .A4(_02260_),
    .ZN(_02261_));
 OAI221_X2 _06499_ (.A(_01350_),
    .B1(_02249_),
    .B2(_02261_),
    .C1(_01064_),
    .C2(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[0][2] ),
    .ZN(_02262_));
 AOI22_X1 _06500_ (.A1(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[25][2] ),
    .A2(net148),
    .B1(net245),
    .B2(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[20][2] ),
    .ZN(_02263_));
 AOI22_X1 _06501_ (.A1(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[16][2] ),
    .A2(net120),
    .B1(net263),
    .B2(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[18][2] ),
    .ZN(_02264_));
 AOI22_X1 _06502_ (.A1(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[26][2] ),
    .A2(net175),
    .B1(net222),
    .B2(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[22][2] ),
    .ZN(_02265_));
 AOI22_X1 _06503_ (.A1(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[23][2] ),
    .A2(net102),
    .B1(net217),
    .B2(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[9][2] ),
    .ZN(_02266_));
 AND4_X1 _06504_ (.A1(_02263_),
    .A2(_02264_),
    .A3(_02265_),
    .A4(_02266_),
    .ZN(_02267_));
 AOI22_X1 _06505_ (.A1(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[24][2] ),
    .A2(net74),
    .B1(net242),
    .B2(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[2][2] ),
    .ZN(_02268_));
 AOI22_X1 _06506_ (.A1(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[7][2] ),
    .A2(_01076_),
    .B1(net126),
    .B2(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[4][2] ),
    .ZN(_02269_));
 MUX2_X1 _06507_ (.A(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[5][2] ),
    .B(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[21][2] ),
    .S(net1),
    .Z(_02270_));
 AOI221_X1 _06508_ (.A(net114),
    .B1(_01597_),
    .B2(_02270_),
    .C1(net158),
    .C2(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[6][2] ),
    .ZN(_02271_));
 NAND4_X1 _06509_ (.A1(_02267_),
    .A2(_02268_),
    .A3(_02269_),
    .A4(_02271_),
    .ZN(_02272_));
 AOI22_X1 _06510_ (.A1(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[15][2] ),
    .A2(net108),
    .B1(net77),
    .B2(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[28][2] ),
    .ZN(_02273_));
 AOI22_X1 _06511_ (.A1(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[8][2] ),
    .A2(net181),
    .B1(net90),
    .B2(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[10][2] ),
    .ZN(_02274_));
 AOI22_X1 _06512_ (.A1(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[12][2] ),
    .A2(net269),
    .B1(net204),
    .B2(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[13][2] ),
    .ZN(_02275_));
 AOI22_X1 _06513_ (.A1(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[17][2] ),
    .A2(net80),
    .B1(net144),
    .B2(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[29][2] ),
    .ZN(_02276_));
 NAND4_X1 _06514_ (.A1(_02273_),
    .A2(_02274_),
    .A3(_02275_),
    .A4(_02276_),
    .ZN(_02277_));
 AOI22_X1 _06515_ (.A1(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[3][2] ),
    .A2(net64),
    .B1(net236),
    .B2(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[11][2] ),
    .ZN(_02278_));
 AOI22_X1 _06516_ (.A1(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[27][2] ),
    .A2(net192),
    .B1(net260),
    .B2(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[1][2] ),
    .ZN(_02279_));
 AOI22_X1 _06517_ (.A1(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[31][2] ),
    .A2(net95),
    .B1(net87),
    .B2(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[14][2] ),
    .ZN(_02280_));
 AOI22_X1 _06518_ (.A1(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[30][2] ),
    .A2(net212),
    .B1(net195),
    .B2(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[19][2] ),
    .ZN(_02281_));
 NAND4_X1 _06519_ (.A1(_02278_),
    .A2(_02279_),
    .A3(_02280_),
    .A4(_02281_),
    .ZN(_02282_));
 NOR3_X1 _06520_ (.A1(_02272_),
    .A2(_02277_),
    .A3(_02282_),
    .ZN(_02283_));
 OAI21_X1 _06521_ (.A(_01700_),
    .B1(net130),
    .B2(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[0][2] ),
    .ZN(_02284_));
 OAI21_X1 _06522_ (.A(_02262_),
    .B1(_02283_),
    .B2(_02284_),
    .ZN(_02285_));
 AOI22_X1 _06523_ (.A1(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[7][2] ),
    .A2(net70),
    .B1(net89),
    .B2(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[10][2] ),
    .ZN(_02286_));
 AOI22_X1 _06524_ (.A1(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[26][2] ),
    .A2(net171),
    .B1(net206),
    .B2(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[13][2] ),
    .ZN(_02287_));
 AOI22_X1 _06525_ (.A1(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[28][2] ),
    .A2(_01032_),
    .B1(net228),
    .B2(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[22][2] ),
    .ZN(_02288_));
 AOI22_X2 _06526_ (.A1(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[29][2] ),
    .A2(net146),
    .B1(net253),
    .B2(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[1][2] ),
    .ZN(_02289_));
 NAND4_X2 _06527_ (.A1(_02286_),
    .A2(_02287_),
    .A3(_02288_),
    .A4(_02289_),
    .ZN(_02290_));
 AOI22_X1 _06528_ (.A1(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[8][2] ),
    .A2(net182),
    .B1(net139),
    .B2(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[5][2] ),
    .ZN(_02291_));
 AOI22_X1 _06529_ (.A1(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[23][2] ),
    .A2(net98),
    .B1(net248),
    .B2(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[20][2] ),
    .ZN(_02292_));
 AOI22_X1 _06530_ (.A1(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[2][2] ),
    .A2(net243),
    .B1(net237),
    .B2(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[11][2] ),
    .ZN(_02293_));
 AOI21_X1 _06531_ (.A(_01119_),
    .B1(net84),
    .B2(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[21][2] ),
    .ZN(_02294_));
 NAND4_X1 _06532_ (.A1(_02291_),
    .A2(_02292_),
    .A3(_02293_),
    .A4(_02294_),
    .ZN(_02295_));
 AOI22_X1 _06533_ (.A1(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[3][2] ),
    .A2(net65),
    .B1(net149),
    .B2(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[25][2] ),
    .ZN(_02296_));
 AOI22_X1 _06534_ (.A1(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[18][2] ),
    .A2(net264),
    .B1(net198),
    .B2(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[19][2] ),
    .ZN(_02297_));
 AOI22_X1 _06535_ (.A1(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[17][2] ),
    .A2(net78),
    .B1(net109),
    .B2(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[15][2] ),
    .ZN(_02298_));
 AOI22_X2 _06536_ (.A1(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[24][2] ),
    .A2(net73),
    .B1(net272),
    .B2(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[12][2] ),
    .ZN(_02299_));
 NAND4_X2 _06537_ (.A1(_02296_),
    .A2(_02297_),
    .A3(_02298_),
    .A4(_02299_),
    .ZN(_02300_));
 TAPCELL_X1 PHY_68 ();
 AOI22_X1 _06539_ (.A1(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[16][2] ),
    .A2(net119),
    .B1(net160),
    .B2(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[6][2] ),
    .ZN(_02302_));
 AOI22_X1 _06540_ (.A1(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[14][2] ),
    .A2(net87),
    .B1(_00999_),
    .B2(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[9][2] ),
    .ZN(_02303_));
 AOI22_X1 _06541_ (.A1(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[31][2] ),
    .A2(_01149_),
    .B1(net128),
    .B2(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[4][2] ),
    .ZN(_02304_));
 AOI22_X1 _06542_ (.A1(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[27][2] ),
    .A2(net192),
    .B1(net211),
    .B2(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[30][2] ),
    .ZN(_02305_));
 NAND4_X1 _06543_ (.A1(_02302_),
    .A2(_02303_),
    .A3(_02304_),
    .A4(_02305_),
    .ZN(_02306_));
 NOR4_X2 _06544_ (.A1(_02290_),
    .A2(_02295_),
    .A3(_02300_),
    .A4(_02306_),
    .ZN(_02307_));
 OAI21_X1 _06545_ (.A(_01408_),
    .B1(net130),
    .B2(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[0][2] ),
    .ZN(_02308_));
 OAI21_X1 _06546_ (.A(_01406_),
    .B1(_02307_),
    .B2(_02308_),
    .ZN(_02309_));
 AOI22_X1 _06547_ (.A1(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[24][2] ),
    .A2(_01059_),
    .B1(_00964_),
    .B2(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[18][2] ),
    .ZN(_02310_));
 AOI22_X1 _06548_ (.A1(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[25][2] ),
    .A2(net147),
    .B1(net141),
    .B2(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[29][2] ),
    .ZN(_02311_));
 AOI22_X1 _06549_ (.A1(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[22][2] ),
    .A2(net227),
    .B1(net203),
    .B2(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[13][2] ),
    .ZN(_02312_));
 TAPCELL_X1 PHY_67 ();
 AOI22_X2 _06551_ (.A1(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[3][2] ),
    .A2(_01102_),
    .B1(_00956_),
    .B2(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[10][2] ),
    .ZN(_02314_));
 NAND4_X2 _06552_ (.A1(_02310_),
    .A2(_02311_),
    .A3(_02312_),
    .A4(_02314_),
    .ZN(_02315_));
 AOI22_X1 _06553_ (.A1(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[12][2] ),
    .A2(net273),
    .B1(net213),
    .B2(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[30][2] ),
    .ZN(_02316_));
 AOI22_X1 _06554_ (.A1(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[28][2] ),
    .A2(net76),
    .B1(net238),
    .B2(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[2][2] ),
    .ZN(_02317_));
 AOI22_X1 _06555_ (.A1(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[4][2] ),
    .A2(net126),
    .B1(net83),
    .B2(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[21][2] ),
    .ZN(_02318_));
 AOI21_X1 _06556_ (.A(net114),
    .B1(net229),
    .B2(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[11][2] ),
    .ZN(_02319_));
 NAND4_X2 _06557_ (.A1(_02316_),
    .A2(_02317_),
    .A3(_02318_),
    .A4(_02319_),
    .ZN(_02320_));
 AOI22_X2 _06558_ (.A1(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[31][2] ),
    .A2(net94),
    .B1(net199),
    .B2(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[19][2] ),
    .ZN(_02321_));
 AOI22_X2 _06559_ (.A1(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[23][2] ),
    .A2(net97),
    .B1(net122),
    .B2(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[16][2] ),
    .ZN(_02322_));
 AOI22_X2 _06560_ (.A1(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[15][2] ),
    .A2(net110),
    .B1(net261),
    .B2(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[1][2] ),
    .ZN(_02323_));
 AOI22_X2 _06561_ (.A1(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[27][2] ),
    .A2(net187),
    .B1(net185),
    .B2(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[8][2] ),
    .ZN(_02324_));
 NAND4_X4 _06562_ (.A1(_02321_),
    .A2(_02322_),
    .A3(_02323_),
    .A4(_02324_),
    .ZN(_02325_));
 AOI22_X1 _06563_ (.A1(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[5][2] ),
    .A2(net133),
    .B1(net88),
    .B2(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[14][2] ),
    .ZN(_02326_));
 TAPCELL_X1 PHY_66 ();
 AOI22_X1 _06565_ (.A1(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[17][2] ),
    .A2(net79),
    .B1(net174),
    .B2(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[26][2] ),
    .ZN(_02328_));
 AOI22_X1 _06566_ (.A1(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[7][2] ),
    .A2(net69),
    .B1(net246),
    .B2(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[20][2] ),
    .ZN(_02329_));
 AOI22_X1 _06567_ (.A1(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[6][2] ),
    .A2(net157),
    .B1(net218),
    .B2(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[9][2] ),
    .ZN(_02330_));
 NAND4_X2 _06568_ (.A1(_02326_),
    .A2(_02328_),
    .A3(_02329_),
    .A4(_02330_),
    .ZN(_02331_));
 NOR4_X4 _06569_ (.A1(_02315_),
    .A2(_02320_),
    .A3(_02325_),
    .A4(_02331_),
    .ZN(_02332_));
 OAI21_X1 _06570_ (.A(_01583_),
    .B1(net130),
    .B2(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[0][2] ),
    .ZN(_02333_));
 AOI22_X1 _06571_ (.A1(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[3][2] ),
    .A2(net63),
    .B1(_01059_),
    .B2(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[24][2] ),
    .ZN(_02334_));
 AOI22_X1 _06572_ (.A1(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[15][2] ),
    .A2(net111),
    .B1(_00989_),
    .B2(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[2][2] ),
    .ZN(_02335_));
 AOI22_X1 _06573_ (.A1(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[14][2] ),
    .A2(net88),
    .B1(net215),
    .B2(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[30][2] ),
    .ZN(_02336_));
 AOI22_X1 _06574_ (.A1(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[16][2] ),
    .A2(net121),
    .B1(net70),
    .B2(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[7][2] ),
    .ZN(_02337_));
 NAND4_X1 _06575_ (.A1(_02334_),
    .A2(_02335_),
    .A3(_02336_),
    .A4(_02337_),
    .ZN(_02338_));
 AOI22_X1 _06576_ (.A1(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[5][2] ),
    .A2(net135),
    .B1(net129),
    .B2(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[4][2] ),
    .ZN(_02339_));
 AOI22_X1 _06577_ (.A1(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[26][2] ),
    .A2(net167),
    .B1(net244),
    .B2(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[20][2] ),
    .ZN(_02340_));
 AOI22_X1 _06578_ (.A1(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[8][2] ),
    .A2(net176),
    .B1(net151),
    .B2(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[25][2] ),
    .ZN(_02341_));
 AOI21_X1 _06579_ (.A(net115),
    .B1(_00996_),
    .B2(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[22][2] ),
    .ZN(_02342_));
 NAND4_X1 _06580_ (.A1(_02339_),
    .A2(_02340_),
    .A3(_02341_),
    .A4(_02342_),
    .ZN(_02343_));
 AOI22_X1 _06581_ (.A1(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[17][2] ),
    .A2(net81),
    .B1(net89),
    .B2(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[10][2] ),
    .ZN(_02344_));
 AOI22_X1 _06582_ (.A1(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[23][2] ),
    .A2(_01144_),
    .B1(_01149_),
    .B2(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[31][2] ),
    .ZN(_02345_));
 AOI22_X1 _06583_ (.A1(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[6][2] ),
    .A2(net156),
    .B1(_00981_),
    .B2(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[21][2] ),
    .ZN(_02346_));
 TAPCELL_X1 PHY_65 ();
 AOI22_X2 _06585_ (.A1(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[27][2] ),
    .A2(net186),
    .B1(_01050_),
    .B2(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[29][2] ),
    .ZN(_02348_));
 NAND4_X2 _06586_ (.A1(_02344_),
    .A2(_02345_),
    .A3(_02346_),
    .A4(_02348_),
    .ZN(_02349_));
 TAPCELL_X1 PHY_64 ();
 AOI22_X1 _06588_ (.A1(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[18][2] ),
    .A2(_00964_),
    .B1(_01007_),
    .B2(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[13][2] ),
    .ZN(_02351_));
 AOI22_X1 _06589_ (.A1(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[12][2] ),
    .A2(net274),
    .B1(net262),
    .B2(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[1][2] ),
    .ZN(_02352_));
 AOI22_X1 _06590_ (.A1(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[9][2] ),
    .A2(net221),
    .B1(net200),
    .B2(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[19][2] ),
    .ZN(_02353_));
 TAPCELL_X1 PHY_63 ();
 AOI22_X2 _06592_ (.A1(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[28][2] ),
    .A2(_01032_),
    .B1(net231),
    .B2(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[11][2] ),
    .ZN(_02355_));
 NAND4_X2 _06593_ (.A1(_02351_),
    .A2(_02352_),
    .A3(_02353_),
    .A4(_02355_),
    .ZN(_02356_));
 NOR4_X2 _06594_ (.A1(_02338_),
    .A2(_02343_),
    .A3(_02349_),
    .A4(_02356_),
    .ZN(_02357_));
 OAI21_X1 _06595_ (.A(_01502_),
    .B1(net130),
    .B2(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[0][2] ),
    .ZN(_02358_));
 OAI22_X2 _06596_ (.A1(_02332_),
    .A2(_02333_),
    .B1(_02357_),
    .B2(_02358_),
    .ZN(_02359_));
 AOI22_X1 _06597_ (.A1(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[27][2] ),
    .A2(net191),
    .B1(net119),
    .B2(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[16][2] ),
    .ZN(_02360_));
 TAPCELL_X1 PHY_62 ();
 AOI22_X1 _06599_ (.A1(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[25][2] ),
    .A2(net149),
    .B1(net207),
    .B2(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[30][2] ),
    .ZN(_02362_));
 AOI22_X1 _06600_ (.A1(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[8][2] ),
    .A2(net182),
    .B1(net84),
    .B2(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[21][2] ),
    .ZN(_02363_));
 TAPCELL_X1 PHY_61 ();
 AOI22_X2 _06602_ (.A1(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[29][2] ),
    .A2(net140),
    .B1(net266),
    .B2(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[12][2] ),
    .ZN(_02365_));
 NAND4_X2 _06603_ (.A1(_02360_),
    .A2(_02362_),
    .A3(_02363_),
    .A4(_02365_),
    .ZN(_02366_));
 AOI22_X1 _06604_ (.A1(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[6][2] ),
    .A2(net160),
    .B1(net223),
    .B2(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[22][2] ),
    .ZN(_02367_));
 AOI22_X1 _06605_ (.A1(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[7][2] ),
    .A2(net67),
    .B1(net87),
    .B2(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[14][2] ),
    .ZN(_02368_));
 AOI21_X1 _06606_ (.A(_01119_),
    .B1(net220),
    .B2(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[9][2] ),
    .ZN(_02369_));
 AOI22_X1 _06607_ (.A1(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[10][2] ),
    .A2(net91),
    .B1(net248),
    .B2(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[20][2] ),
    .ZN(_02370_));
 NAND4_X1 _06608_ (.A1(_02367_),
    .A2(_02368_),
    .A3(_02369_),
    .A4(_02370_),
    .ZN(_02371_));
 AOI22_X1 _06609_ (.A1(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[28][2] ),
    .A2(net75),
    .B1(net232),
    .B2(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[11][2] ),
    .ZN(_02372_));
 AOI22_X1 _06610_ (.A1(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[23][2] ),
    .A2(net98),
    .B1(_01149_),
    .B2(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[31][2] ),
    .ZN(_02373_));
 AOI22_X1 _06611_ (.A1(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[24][2] ),
    .A2(net72),
    .B1(net206),
    .B2(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[13][2] ),
    .ZN(_02374_));
 AOI22_X1 _06612_ (.A1(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[26][2] ),
    .A2(net168),
    .B1(net198),
    .B2(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[19][2] ),
    .ZN(_02375_));
 NAND4_X1 _06613_ (.A1(_02372_),
    .A2(_02373_),
    .A3(_02374_),
    .A4(_02375_),
    .ZN(_02376_));
 AOI22_X1 _06614_ (.A1(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[5][2] ),
    .A2(net136),
    .B1(net243),
    .B2(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[2][2] ),
    .ZN(_02377_));
 TAPCELL_X1 PHY_60 ();
 AOI22_X1 _06616_ (.A1(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[15][2] ),
    .A2(net109),
    .B1(net264),
    .B2(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[18][2] ),
    .ZN(_02379_));
 AOI22_X1 _06617_ (.A1(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[4][2] ),
    .A2(net128),
    .B1(net258),
    .B2(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[1][2] ),
    .ZN(_02380_));
 AOI22_X2 _06618_ (.A1(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[17][2] ),
    .A2(net78),
    .B1(net65),
    .B2(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[3][2] ),
    .ZN(_02381_));
 NAND4_X2 _06619_ (.A1(_02377_),
    .A2(_02379_),
    .A3(_02380_),
    .A4(_02381_),
    .ZN(_02382_));
 NOR4_X2 _06620_ (.A1(_02366_),
    .A2(_02371_),
    .A3(_02376_),
    .A4(_02382_),
    .ZN(_02383_));
 OAI21_X1 _06621_ (.A(_00923_),
    .B1(_01064_),
    .B2(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[0][2] ),
    .ZN(_02384_));
 AOI22_X1 _06622_ (.A1(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[28][2] ),
    .A2(net75),
    .B1(net72),
    .B2(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[24][2] ),
    .ZN(_02385_));
 AOI22_X1 _06623_ (.A1(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[2][2] ),
    .A2(net243),
    .B1(net220),
    .B2(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[9][2] ),
    .ZN(_02386_));
 AOI22_X1 _06624_ (.A1(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[26][2] ),
    .A2(net168),
    .B1(net197),
    .B2(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[19][2] ),
    .ZN(_02387_));
 AOI22_X1 _06625_ (.A1(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[3][2] ),
    .A2(net65),
    .B1(net118),
    .B2(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[16][2] ),
    .ZN(_02388_));
 NAND4_X1 _06626_ (.A1(_02385_),
    .A2(_02386_),
    .A3(_02387_),
    .A4(_02388_),
    .ZN(_02389_));
 AOI22_X1 _06627_ (.A1(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[8][2] ),
    .A2(net183),
    .B1(net82),
    .B2(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[21][2] ),
    .ZN(_02390_));
 AOI22_X1 _06628_ (.A1(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[27][2] ),
    .A2(net189),
    .B1(net86),
    .B2(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[14][2] ),
    .ZN(_02391_));
 AOI22_X1 _06629_ (.A1(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[18][2] ),
    .A2(net264),
    .B1(net232),
    .B2(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[11][2] ),
    .ZN(_02392_));
 AOI21_X1 _06630_ (.A(_01119_),
    .B1(net207),
    .B2(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[30][2] ),
    .ZN(_02393_));
 NAND4_X2 _06631_ (.A1(_02390_),
    .A2(_02391_),
    .A3(_02392_),
    .A4(_02393_),
    .ZN(_02394_));
 AOI22_X1 _06632_ (.A1(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[25][2] ),
    .A2(net149),
    .B1(net136),
    .B2(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[5][2] ),
    .ZN(_02395_));
 AOI22_X1 _06633_ (.A1(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[17][2] ),
    .A2(net78),
    .B1(net96),
    .B2(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[31][2] ),
    .ZN(_02396_));
 TAPCELL_X1 PHY_59 ();
 AOI22_X1 _06635_ (.A1(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[29][2] ),
    .A2(net140),
    .B1(net266),
    .B2(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[12][2] ),
    .ZN(_02398_));
 AOI22_X2 _06636_ (.A1(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[22][2] ),
    .A2(net223),
    .B1(net206),
    .B2(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[13][2] ),
    .ZN(_02399_));
 NAND4_X2 _06637_ (.A1(_02395_),
    .A2(_02396_),
    .A3(_02398_),
    .A4(_02399_),
    .ZN(_02400_));
 AOI22_X1 _06638_ (.A1(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[4][2] ),
    .A2(net125),
    .B1(net91),
    .B2(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[10][2] ),
    .ZN(_02401_));
 AOI22_X1 _06639_ (.A1(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[23][2] ),
    .A2(net103),
    .B1(net161),
    .B2(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[6][2] ),
    .ZN(_02402_));
 AOI22_X1 _06640_ (.A1(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[7][2] ),
    .A2(net67),
    .B1(net247),
    .B2(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[20][2] ),
    .ZN(_02403_));
 AOI22_X2 _06641_ (.A1(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[15][2] ),
    .A2(net106),
    .B1(net257),
    .B2(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[1][2] ),
    .ZN(_02404_));
 NAND4_X2 _06642_ (.A1(_02401_),
    .A2(_02402_),
    .A3(_02403_),
    .A4(_02404_),
    .ZN(_02405_));
 NOR4_X2 _06643_ (.A1(_02389_),
    .A2(_02394_),
    .A3(_02400_),
    .A4(_02405_),
    .ZN(_02406_));
 OAI21_X1 _06644_ (.A(_01164_),
    .B1(_01064_),
    .B2(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[0][2] ),
    .ZN(_02407_));
 OAI22_X2 _06645_ (.A1(_02383_),
    .A2(_02384_),
    .B1(_02406_),
    .B2(_02407_),
    .ZN(_02408_));
 NOR4_X2 _06646_ (.A1(_02285_),
    .A2(_02309_),
    .A3(_02359_),
    .A4(_02408_),
    .ZN(_02409_));
 AOI22_X1 _06647_ (.A1(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[21][2] ),
    .A2(_00981_),
    .B1(net231),
    .B2(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[11][2] ),
    .ZN(_02410_));
 AOI22_X1 _06648_ (.A1(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[15][2] ),
    .A2(net112),
    .B1(net274),
    .B2(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[12][2] ),
    .ZN(_02411_));
 TAPCELL_X1 PHY_58 ();
 AOI22_X1 _06650_ (.A1(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[8][2] ),
    .A2(net176),
    .B1(_00971_),
    .B2(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[14][2] ),
    .ZN(_02413_));
 AOI22_X2 _06651_ (.A1(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[28][2] ),
    .A2(_01032_),
    .B1(net73),
    .B2(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[24][2] ),
    .ZN(_02414_));
 NAND4_X2 _06652_ (.A1(_02410_),
    .A2(_02411_),
    .A3(_02413_),
    .A4(_02414_),
    .ZN(_02415_));
 AOI22_X1 _06653_ (.A1(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[25][2] ),
    .A2(net150),
    .B1(net206),
    .B2(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[13][2] ),
    .ZN(_02416_));
 AOI22_X1 _06654_ (.A1(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[6][2] ),
    .A2(net156),
    .B1(net244),
    .B2(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[20][2] ),
    .ZN(_02417_));
 AOI22_X1 _06655_ (.A1(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[7][2] ),
    .A2(net70),
    .B1(net215),
    .B2(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[30][2] ),
    .ZN(_02418_));
 AOI21_X1 _06656_ (.A(net115),
    .B1(net146),
    .B2(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[29][2] ),
    .ZN(_02419_));
 NAND4_X2 _06657_ (.A1(_02416_),
    .A2(_02417_),
    .A3(_02418_),
    .A4(_02419_),
    .ZN(_02420_));
 AOI22_X1 _06658_ (.A1(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[3][2] ),
    .A2(net63),
    .B1(net228),
    .B2(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[22][2] ),
    .ZN(_02421_));
 AOI22_X1 _06659_ (.A1(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[27][2] ),
    .A2(net186),
    .B1(_00999_),
    .B2(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[9][2] ),
    .ZN(_02422_));
 AOI22_X1 _06660_ (.A1(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[26][2] ),
    .A2(net171),
    .B1(net264),
    .B2(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[18][2] ),
    .ZN(_02423_));
 AOI22_X2 _06661_ (.A1(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[17][2] ),
    .A2(net81),
    .B1(_00989_),
    .B2(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[2][2] ),
    .ZN(_02424_));
 NAND4_X2 _06662_ (.A1(_02421_),
    .A2(_02422_),
    .A3(_02423_),
    .A4(_02424_),
    .ZN(_02425_));
 AOI22_X1 _06663_ (.A1(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[4][2] ),
    .A2(net128),
    .B1(net89),
    .B2(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[10][2] ),
    .ZN(_02426_));
 AOI22_X1 _06664_ (.A1(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[23][2] ),
    .A2(net99),
    .B1(net121),
    .B2(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[16][2] ),
    .ZN(_02427_));
 TAPCELL_X1 PHY_57 ();
 AOI22_X1 _06666_ (.A1(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[31][2] ),
    .A2(_01149_),
    .B1(net253),
    .B2(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[1][2] ),
    .ZN(_02429_));
 AOI22_X2 _06667_ (.A1(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[5][2] ),
    .A2(net135),
    .B1(net201),
    .B2(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[19][2] ),
    .ZN(_02430_));
 NAND4_X2 _06668_ (.A1(_02426_),
    .A2(_02427_),
    .A3(_02429_),
    .A4(_02430_),
    .ZN(_02431_));
 NOR4_X4 _06669_ (.A1(_02415_),
    .A2(_02420_),
    .A3(_02425_),
    .A4(_02431_),
    .ZN(_02432_));
 OAI21_X1 _06670_ (.A(_01731_),
    .B1(net130),
    .B2(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[0][2] ),
    .ZN(_02433_));
 AOI22_X1 _06671_ (.A1(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[28][2] ),
    .A2(net77),
    .B1(net204),
    .B2(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[13][2] ),
    .ZN(_02434_));
 AOI22_X1 _06672_ (.A1(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[8][2] ),
    .A2(net179),
    .B1(net242),
    .B2(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[2][2] ),
    .ZN(_02435_));
 AOI22_X1 _06673_ (.A1(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[11][2] ),
    .A2(net234),
    .B1(net219),
    .B2(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[9][2] ),
    .ZN(_02436_));
 AOI22_X1 _06674_ (.A1(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[5][2] ),
    .A2(net132),
    .B1(net68),
    .B2(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[7][2] ),
    .ZN(_02437_));
 NAND4_X1 _06675_ (.A1(_02434_),
    .A2(_02435_),
    .A3(_02436_),
    .A4(_02437_),
    .ZN(_02438_));
 AOI22_X1 _06676_ (.A1(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[17][2] ),
    .A2(net80),
    .B1(net224),
    .B2(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[22][2] ),
    .ZN(_02439_));
 AOI22_X1 _06677_ (.A1(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[3][2] ),
    .A2(net64),
    .B1(net153),
    .B2(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[25][2] ),
    .ZN(_02440_));
 AOI22_X1 _06678_ (.A1(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[31][2] ),
    .A2(net95),
    .B1(net82),
    .B2(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[21][2] ),
    .ZN(_02441_));
 AOI21_X1 _06679_ (.A(net113),
    .B1(net256),
    .B2(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[1][2] ),
    .ZN(_02442_));
 NAND4_X1 _06680_ (.A1(_02439_),
    .A2(_02440_),
    .A3(_02441_),
    .A4(_02442_),
    .ZN(_02443_));
 AOI22_X1 _06681_ (.A1(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[15][2] ),
    .A2(net106),
    .B1(net74),
    .B2(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[24][2] ),
    .ZN(_02444_));
 AOI22_X1 _06682_ (.A1(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[27][2] ),
    .A2(net190),
    .B1(net265),
    .B2(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[18][2] ),
    .ZN(_02445_));
 AOI22_X1 _06683_ (.A1(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[16][2] ),
    .A2(net117),
    .B1(net90),
    .B2(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[10][2] ),
    .ZN(_02446_));
 AOI22_X1 _06684_ (.A1(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[23][2] ),
    .A2(net101),
    .B1(net163),
    .B2(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[6][2] ),
    .ZN(_02447_));
 NAND4_X1 _06685_ (.A1(_02444_),
    .A2(_02445_),
    .A3(_02446_),
    .A4(_02447_),
    .ZN(_02448_));
 AOI22_X1 _06686_ (.A1(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[14][2] ),
    .A2(net85),
    .B1(net251),
    .B2(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[20][2] ),
    .ZN(_02449_));
 AOI22_X1 _06687_ (.A1(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[12][2] ),
    .A2(net269),
    .B1(net194),
    .B2(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[19][2] ),
    .ZN(_02450_));
 AOI22_X1 _06688_ (.A1(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[4][2] ),
    .A2(net124),
    .B1(net209),
    .B2(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[30][2] ),
    .ZN(_02451_));
 AOI22_X1 _06689_ (.A1(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[26][2] ),
    .A2(net170),
    .B1(net142),
    .B2(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[29][2] ),
    .ZN(_02452_));
 NAND4_X1 _06690_ (.A1(_02449_),
    .A2(_02450_),
    .A3(_02451_),
    .A4(_02452_),
    .ZN(_02453_));
 NOR4_X2 _06691_ (.A1(_02438_),
    .A2(_02443_),
    .A3(_02448_),
    .A4(_02453_),
    .ZN(_02454_));
 OAI21_X1 _06692_ (.A(_01539_),
    .B1(net130),
    .B2(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[0][2] ),
    .ZN(_02455_));
 OAI22_X1 _06693_ (.A1(_02432_),
    .A2(_02433_),
    .B1(_02454_),
    .B2(_02455_),
    .ZN(_02456_));
 AOI22_X1 _06694_ (.A1(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[4][2] ),
    .A2(net123),
    .B1(net193),
    .B2(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[19][2] ),
    .ZN(_02457_));
 AOI22_X1 _06695_ (.A1(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[16][2] ),
    .A2(net116),
    .B1(net87),
    .B2(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[14][2] ),
    .ZN(_02458_));
 AOI22_X1 _06696_ (.A1(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[2][2] ),
    .A2(net240),
    .B1(net208),
    .B2(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[30][2] ),
    .ZN(_02459_));
 AOI22_X1 _06697_ (.A1(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[3][2] ),
    .A2(net66),
    .B1(net83),
    .B2(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[21][2] ),
    .ZN(_02460_));
 NAND4_X1 _06698_ (.A1(_02457_),
    .A2(_02458_),
    .A3(_02459_),
    .A4(_02460_),
    .ZN(_02461_));
 AOI22_X1 _06699_ (.A1(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[26][2] ),
    .A2(net173),
    .B1(net217),
    .B2(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[9][2] ),
    .ZN(_02462_));
 AOI22_X1 _06700_ (.A1(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[17][2] ),
    .A2(net79),
    .B1(net131),
    .B2(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[5][2] ),
    .ZN(_02463_));
 AOI22_X1 _06701_ (.A1(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[24][2] ),
    .A2(net71),
    .B1(net68),
    .B2(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[7][2] ),
    .ZN(_02464_));
 AOI21_X1 _06702_ (.A(net114),
    .B1(net107),
    .B2(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[15][2] ),
    .ZN(_02465_));
 NAND4_X2 _06703_ (.A1(_02462_),
    .A2(_02463_),
    .A3(_02464_),
    .A4(_02465_),
    .ZN(_02466_));
 AOI22_X1 _06704_ (.A1(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[28][2] ),
    .A2(net76),
    .B1(net250),
    .B2(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[20][2] ),
    .ZN(_02467_));
 AOI22_X1 _06705_ (.A1(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[29][2] ),
    .A2(net144),
    .B1(net222),
    .B2(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[22][2] ),
    .ZN(_02468_));
 AOI22_X1 _06706_ (.A1(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[27][2] ),
    .A2(net188),
    .B1(net93),
    .B2(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[31][2] ),
    .ZN(_02469_));
 AOI22_X2 _06707_ (.A1(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[23][2] ),
    .A2(net100),
    .B1(net90),
    .B2(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[10][2] ),
    .ZN(_02470_));
 NAND4_X2 _06708_ (.A1(_02467_),
    .A2(_02468_),
    .A3(_02469_),
    .A4(_02470_),
    .ZN(_02471_));
 AOI22_X1 _06709_ (.A1(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[25][2] ),
    .A2(net152),
    .B1(net268),
    .B2(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[12][2] ),
    .ZN(_02472_));
 AOI22_X1 _06710_ (.A1(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[1][2] ),
    .A2(net254),
    .B1(net236),
    .B2(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[11][2] ),
    .ZN(_02473_));
 AOI22_X1 _06711_ (.A1(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[18][2] ),
    .A2(net263),
    .B1(net204),
    .B2(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[13][2] ),
    .ZN(_02474_));
 AOI22_X1 _06712_ (.A1(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[8][2] ),
    .A2(net180),
    .B1(net162),
    .B2(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[6][2] ),
    .ZN(_02475_));
 NAND4_X1 _06713_ (.A1(_02472_),
    .A2(_02473_),
    .A3(_02474_),
    .A4(_02475_),
    .ZN(_02476_));
 NOR4_X2 _06714_ (.A1(_02461_),
    .A2(_02466_),
    .A3(_02471_),
    .A4(_02476_),
    .ZN(_02477_));
 OAI21_X1 _06715_ (.A(_01401_),
    .B1(net130),
    .B2(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[0][2] ),
    .ZN(_02478_));
 AOI22_X1 _06716_ (.A1(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[31][2] ),
    .A2(net94),
    .B1(_01007_),
    .B2(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[13][2] ),
    .ZN(_02479_));
 AOI22_X1 _06717_ (.A1(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[16][2] ),
    .A2(net122),
    .B1(net221),
    .B2(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[9][2] ),
    .ZN(_02480_));
 AOI22_X1 _06718_ (.A1(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[6][2] ),
    .A2(net159),
    .B1(_00993_),
    .B2(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[11][2] ),
    .ZN(_02481_));
 AOI22_X1 _06719_ (.A1(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[27][2] ),
    .A2(net186),
    .B1(net239),
    .B2(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[2][2] ),
    .ZN(_02482_));
 NAND4_X2 _06720_ (.A1(_02479_),
    .A2(_02480_),
    .A3(_02481_),
    .A4(_02482_),
    .ZN(_02483_));
 AOI22_X1 _06721_ (.A1(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[14][2] ),
    .A2(net88),
    .B1(net200),
    .B2(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[19][2] ),
    .ZN(_02484_));
 AOI22_X1 _06722_ (.A1(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[3][2] ),
    .A2(net63),
    .B1(net216),
    .B2(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[30][2] ),
    .ZN(_02485_));
 MUX2_X1 _06723_ (.A(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[5][2] ),
    .B(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[21][2] ),
    .S(net1),
    .Z(_02486_));
 AOI221_X1 _06724_ (.A(net115),
    .B1(_01597_),
    .B2(_02486_),
    .C1(net246),
    .C2(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[20][2] ),
    .ZN(_02487_));
 NAND3_X1 _06725_ (.A1(_02484_),
    .A2(_02485_),
    .A3(_02487_),
    .ZN(_02488_));
 AOI22_X1 _06726_ (.A1(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[23][2] ),
    .A2(net97),
    .B1(net89),
    .B2(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[10][2] ),
    .ZN(_02489_));
 AOI22_X1 _06727_ (.A1(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[26][2] ),
    .A2(net167),
    .B1(net262),
    .B2(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[1][2] ),
    .ZN(_02490_));
 AOI22_X1 _06728_ (.A1(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[28][2] ),
    .A2(net76),
    .B1(net129),
    .B2(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[4][2] ),
    .ZN(_02491_));
 AOI22_X2 _06729_ (.A1(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[18][2] ),
    .A2(_00964_),
    .B1(net227),
    .B2(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[22][2] ),
    .ZN(_02492_));
 NAND4_X2 _06730_ (.A1(_02489_),
    .A2(_02490_),
    .A3(_02491_),
    .A4(_02492_),
    .ZN(_02493_));
 AOI22_X1 _06731_ (.A1(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[25][2] ),
    .A2(net151),
    .B1(net273),
    .B2(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[12][2] ),
    .ZN(_02494_));
 AOI22_X1 _06732_ (.A1(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[17][2] ),
    .A2(net81),
    .B1(net141),
    .B2(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[29][2] ),
    .ZN(_02495_));
 AOI22_X1 _06733_ (.A1(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[24][2] ),
    .A2(_01059_),
    .B1(net70),
    .B2(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[7][2] ),
    .ZN(_02496_));
 AOI22_X1 _06734_ (.A1(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[15][2] ),
    .A2(net110),
    .B1(net185),
    .B2(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[8][2] ),
    .ZN(_02497_));
 NAND4_X1 _06735_ (.A1(_02494_),
    .A2(_02495_),
    .A3(_02496_),
    .A4(_02497_),
    .ZN(_02498_));
 NOR4_X2 _06736_ (.A1(_02483_),
    .A2(_02488_),
    .A3(_02493_),
    .A4(_02498_),
    .ZN(_02499_));
 OAI21_X1 _06737_ (.A(_01662_),
    .B1(net130),
    .B2(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[0][2] ),
    .ZN(_02500_));
 OAI22_X1 _06738_ (.A1(_02477_),
    .A2(_02478_),
    .B1(_02499_),
    .B2(_02500_),
    .ZN(_02501_));
 AOI22_X1 _06739_ (.A1(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[5][2] ),
    .A2(net133),
    .B1(_00964_),
    .B2(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[18][2] ),
    .ZN(_02502_));
 AOI22_X1 _06740_ (.A1(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[26][2] ),
    .A2(net166),
    .B1(net246),
    .B2(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[20][2] ),
    .ZN(_02503_));
 AOI22_X1 _06741_ (.A1(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[12][2] ),
    .A2(net273),
    .B1(net214),
    .B2(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[30][2] ),
    .ZN(_02504_));
 AOI22_X1 _06742_ (.A1(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[17][2] ),
    .A2(net81),
    .B1(net239),
    .B2(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[2][2] ),
    .ZN(_02505_));
 NAND4_X1 _06743_ (.A1(_02502_),
    .A2(_02503_),
    .A3(_02504_),
    .A4(_02505_),
    .ZN(_02506_));
 AOI22_X1 _06744_ (.A1(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[6][2] ),
    .A2(net159),
    .B1(net88),
    .B2(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[14][2] ),
    .ZN(_02507_));
 AOI22_X1 _06745_ (.A1(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[4][2] ),
    .A2(net127),
    .B1(net218),
    .B2(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[9][2] ),
    .ZN(_02508_));
 AOI22_X1 _06746_ (.A1(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[10][2] ),
    .A2(net89),
    .B1(net203),
    .B2(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[13][2] ),
    .ZN(_02509_));
 AOI21_X1 _06747_ (.A(net115),
    .B1(net261),
    .B2(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[1][2] ),
    .ZN(_02510_));
 NAND4_X2 _06748_ (.A1(_02507_),
    .A2(_02508_),
    .A3(_02509_),
    .A4(_02510_),
    .ZN(_02511_));
 AOI22_X1 _06749_ (.A1(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[27][2] ),
    .A2(net187),
    .B1(net227),
    .B2(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[22][2] ),
    .ZN(_02512_));
 AOI22_X1 _06750_ (.A1(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[25][2] ),
    .A2(net147),
    .B1(_01059_),
    .B2(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[24][2] ),
    .ZN(_02513_));
 AOI22_X1 _06751_ (.A1(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[29][2] ),
    .A2(net141),
    .B1(_00981_),
    .B2(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[21][2] ),
    .ZN(_02514_));
 AOI22_X1 _06752_ (.A1(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[11][2] ),
    .A2(net230),
    .B1(net202),
    .B2(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[19][2] ),
    .ZN(_02515_));
 NAND4_X1 _06753_ (.A1(_02512_),
    .A2(_02513_),
    .A3(_02514_),
    .A4(_02515_),
    .ZN(_02516_));
 AOI22_X1 _06754_ (.A1(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[23][2] ),
    .A2(net97),
    .B1(net110),
    .B2(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[15][2] ),
    .ZN(_02517_));
 AOI22_X2 _06755_ (.A1(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[16][2] ),
    .A2(net122),
    .B1(net177),
    .B2(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[8][2] ),
    .ZN(_02518_));
 AOI22_X1 _06756_ (.A1(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[3][2] ),
    .A2(net63),
    .B1(net76),
    .B2(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[28][2] ),
    .ZN(_02519_));
 AOI22_X2 _06757_ (.A1(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[7][2] ),
    .A2(net70),
    .B1(net94),
    .B2(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[31][2] ),
    .ZN(_02520_));
 NAND4_X2 _06758_ (.A1(_02517_),
    .A2(_02518_),
    .A3(_02519_),
    .A4(_02520_),
    .ZN(_02521_));
 NOR4_X2 _06759_ (.A1(_02506_),
    .A2(_02511_),
    .A3(_02516_),
    .A4(_02521_),
    .ZN(_02522_));
 OAI21_X1 _06760_ (.A(_01623_),
    .B1(net130),
    .B2(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[0][2] ),
    .ZN(_02523_));
 AOI22_X1 _06761_ (.A1(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[1][2] ),
    .A2(net254),
    .B1(net83),
    .B2(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[21][2] ),
    .ZN(_02524_));
 AOI22_X1 _06762_ (.A1(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[6][2] ),
    .A2(net158),
    .B1(net240),
    .B2(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[2][2] ),
    .ZN(_02525_));
 AOI22_X1 _06763_ (.A1(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[18][2] ),
    .A2(net263),
    .B1(net87),
    .B2(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[14][2] ),
    .ZN(_02526_));
 AOI22_X1 _06764_ (.A1(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[31][2] ),
    .A2(net93),
    .B1(net268),
    .B2(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[12][2] ),
    .ZN(_02527_));
 NAND4_X1 _06765_ (.A1(_02524_),
    .A2(_02525_),
    .A3(_02526_),
    .A4(_02527_),
    .ZN(_02528_));
 AOI22_X1 _06766_ (.A1(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[17][2] ),
    .A2(net79),
    .B1(net102),
    .B2(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[23][2] ),
    .ZN(_02529_));
 AOI22_X1 _06767_ (.A1(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[10][2] ),
    .A2(_00956_),
    .B1(net213),
    .B2(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[30][2] ),
    .ZN(_02530_));
 AOI22_X1 _06768_ (.A1(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[5][2] ),
    .A2(net134),
    .B1(net222),
    .B2(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[22][2] ),
    .ZN(_02531_));
 AOI21_X1 _06769_ (.A(net114),
    .B1(net120),
    .B2(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[16][2] ),
    .ZN(_02532_));
 NAND4_X1 _06770_ (.A1(_02529_),
    .A2(_02530_),
    .A3(_02531_),
    .A4(_02532_),
    .ZN(_02533_));
 AOI22_X1 _06771_ (.A1(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[25][2] ),
    .A2(net152),
    .B1(net144),
    .B2(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[29][2] ),
    .ZN(_02534_));
 AOI22_X1 _06772_ (.A1(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[3][2] ),
    .A2(net66),
    .B1(net245),
    .B2(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[20][2] ),
    .ZN(_02535_));
 AOI22_X1 _06773_ (.A1(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[8][2] ),
    .A2(net178),
    .B1(net174),
    .B2(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[26][2] ),
    .ZN(_02536_));
 AOI22_X1 _06774_ (.A1(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[15][2] ),
    .A2(net108),
    .B1(net71),
    .B2(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[24][2] ),
    .ZN(_02537_));
 NAND4_X2 _06775_ (.A1(_02534_),
    .A2(_02535_),
    .A3(_02536_),
    .A4(_02537_),
    .ZN(_02538_));
 AOI22_X1 _06776_ (.A1(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[4][2] ),
    .A2(net126),
    .B1(net203),
    .B2(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[13][2] ),
    .ZN(_02539_));
 AOI22_X1 _06777_ (.A1(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[27][2] ),
    .A2(net188),
    .B1(net196),
    .B2(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[19][2] ),
    .ZN(_02540_));
 AOI22_X1 _06778_ (.A1(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[11][2] ),
    .A2(net229),
    .B1(net218),
    .B2(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[9][2] ),
    .ZN(_02541_));
 AOI22_X2 _06779_ (.A1(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[28][2] ),
    .A2(net76),
    .B1(net69),
    .B2(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[7][2] ),
    .ZN(_02542_));
 NAND4_X2 _06780_ (.A1(_02539_),
    .A2(_02540_),
    .A3(_02541_),
    .A4(_02542_),
    .ZN(_02543_));
 NOR4_X2 _06781_ (.A1(_02528_),
    .A2(_02533_),
    .A3(_02538_),
    .A4(_02543_),
    .ZN(_02544_));
 OAI21_X1 _06782_ (.A(_01295_),
    .B1(net130),
    .B2(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[0][2] ),
    .ZN(_02545_));
 OAI22_X2 _06783_ (.A1(_02522_),
    .A2(_02523_),
    .B1(_02544_),
    .B2(_02545_),
    .ZN(_02546_));
 AOI22_X1 _06784_ (.A1(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[8][2] ),
    .A2(_01034_),
    .B1(_01009_),
    .B2(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[19][2] ),
    .ZN(_02547_));
 AOI22_X1 _06785_ (.A1(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[5][2] ),
    .A2(net139),
    .B1(net242),
    .B2(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[2][2] ),
    .ZN(_02548_));
 AND2_X1 _06786_ (.A1(_02547_),
    .A2(_02548_),
    .ZN(_02549_));
 INV_X1 _06787_ (.A(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[31][2] ),
    .ZN(_02550_));
 INV_X1 _06788_ (.A(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[20][2] ),
    .ZN(_02551_));
 OAI22_X1 _06789_ (.A1(_02550_),
    .A2(_00934_),
    .B1(_01691_),
    .B2(_02551_),
    .ZN(_02552_));
 AOI221_X1 _06790_ (.A(_02552_),
    .B1(_01076_),
    .B2(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[7][2] ),
    .C1(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[28][2] ),
    .C2(net77),
    .ZN(_02553_));
 INV_X1 _06791_ (.A(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[27][2] ),
    .ZN(_02554_));
 NAND3_X4 _06792_ (.A1(_00946_),
    .A2(_00926_),
    .A3(_01418_),
    .ZN(_02555_));
 NAND4_X4 _06793_ (.A1(_00911_),
    .A2(net8),
    .A3(_00946_),
    .A4(_01418_),
    .ZN(_02556_));
 INV_X1 _06794_ (.A(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[11][2] ),
    .ZN(_02557_));
 OAI22_X1 _06795_ (.A1(_02554_),
    .A2(_02555_),
    .B1(_02556_),
    .B2(_02557_),
    .ZN(_02558_));
 AOI221_X1 _06796_ (.A(_02558_),
    .B1(net78),
    .B2(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[17][2] ),
    .C1(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[25][2] ),
    .C2(_01046_),
    .ZN(_02559_));
 INV_X1 _06797_ (.A(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[6][2] ),
    .ZN(_02560_));
 OAI21_X1 _06798_ (.A(_01064_),
    .B1(_01681_),
    .B2(_02560_),
    .ZN(_02561_));
 AOI221_X1 _06799_ (.A(_02561_),
    .B1(net65),
    .B2(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[3][2] ),
    .C1(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[24][2] ),
    .C2(net73),
    .ZN(_02562_));
 AND4_X1 _06800_ (.A1(_02549_),
    .A2(_02553_),
    .A3(_02559_),
    .A4(_02562_),
    .ZN(_02563_));
 AOI22_X1 _06801_ (.A1(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[29][2] ),
    .A2(net143),
    .B1(net259),
    .B2(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[1][2] ),
    .ZN(_02564_));
 AOI22_X1 _06802_ (.A1(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[26][2] ),
    .A2(net169),
    .B1(net86),
    .B2(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[14][2] ),
    .ZN(_02565_));
 AOI22_X1 _06803_ (.A1(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[15][2] ),
    .A2(_01123_),
    .B1(net205),
    .B2(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[13][2] ),
    .ZN(_02566_));
 AOI22_X1 _06804_ (.A1(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[9][2] ),
    .A2(net220),
    .B1(net211),
    .B2(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[30][2] ),
    .ZN(_02567_));
 AND4_X1 _06805_ (.A1(_02564_),
    .A2(_02565_),
    .A3(_02566_),
    .A4(_02567_),
    .ZN(_02568_));
 AOI22_X1 _06806_ (.A1(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[23][2] ),
    .A2(net105),
    .B1(net125),
    .B2(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[4][2] ),
    .ZN(_02569_));
 AOI22_X1 _06807_ (.A1(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[16][2] ),
    .A2(net118),
    .B1(net91),
    .B2(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[10][2] ),
    .ZN(_02570_));
 AND2_X1 _06808_ (.A1(_02569_),
    .A2(_02570_),
    .ZN(_02571_));
 AOI22_X1 _06809_ (.A1(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[21][2] ),
    .A2(net83),
    .B1(net224),
    .B2(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[22][2] ),
    .ZN(_02572_));
 AOI22_X1 _06810_ (.A1(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[12][2] ),
    .A2(net271),
    .B1(net265),
    .B2(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[18][2] ),
    .ZN(_02573_));
 AND2_X1 _06811_ (.A1(_02572_),
    .A2(_02573_),
    .ZN(_02574_));
 AND4_X1 _06812_ (.A1(_02563_),
    .A2(_02568_),
    .A3(_02571_),
    .A4(_02574_),
    .ZN(_02575_));
 OAI21_X1 _06813_ (.A(_01764_),
    .B1(net130),
    .B2(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[0][2] ),
    .ZN(_02576_));
 AOI22_X1 _06814_ (.A1(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[4][2] ),
    .A2(net124),
    .B1(net270),
    .B2(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[12][2] ),
    .ZN(_02577_));
 AOI22_X1 _06815_ (.A1(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[5][2] ),
    .A2(net137),
    .B1(net82),
    .B2(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[21][2] ),
    .ZN(_02578_));
 AOI22_X1 _06816_ (.A1(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[24][2] ),
    .A2(net74),
    .B1(net85),
    .B2(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[14][2] ),
    .ZN(_02579_));
 AOI22_X1 _06817_ (.A1(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[8][2] ),
    .A2(net184),
    .B1(net210),
    .B2(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[30][2] ),
    .ZN(_02580_));
 NAND4_X1 _06818_ (.A1(_02577_),
    .A2(_02578_),
    .A3(_02579_),
    .A4(_02580_),
    .ZN(_02581_));
 AOI22_X1 _06819_ (.A1(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[27][2] ),
    .A2(net189),
    .B1(net205),
    .B2(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[13][2] ),
    .ZN(_02582_));
 AOI22_X1 _06820_ (.A1(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[9][2] ),
    .A2(net219),
    .B1(net195),
    .B2(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[19][2] ),
    .ZN(_02583_));
 AOI22_X1 _06821_ (.A1(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[25][2] ),
    .A2(net154),
    .B1(net67),
    .B2(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[7][2] ),
    .ZN(_02584_));
 AOI21_X1 _06822_ (.A(net113),
    .B1(net96),
    .B2(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[31][2] ),
    .ZN(_02585_));
 NAND4_X1 _06823_ (.A1(_02582_),
    .A2(_02583_),
    .A3(_02584_),
    .A4(_02585_),
    .ZN(_02586_));
 AOI22_X1 _06824_ (.A1(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[3][2] ),
    .A2(net64),
    .B1(net163),
    .B2(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[6][2] ),
    .ZN(_02587_));
 AOI22_X1 _06825_ (.A1(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[17][2] ),
    .A2(net80),
    .B1(net234),
    .B2(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[11][2] ),
    .ZN(_02588_));
 AOI22_X1 _06826_ (.A1(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[10][2] ),
    .A2(net90),
    .B1(net247),
    .B2(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[20][2] ),
    .ZN(_02589_));
 AOI22_X2 _06827_ (.A1(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[28][2] ),
    .A2(net75),
    .B1(net265),
    .B2(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[18][2] ),
    .ZN(_02590_));
 NAND4_X2 _06828_ (.A1(_02587_),
    .A2(_02588_),
    .A3(_02589_),
    .A4(_02590_),
    .ZN(_02591_));
 AOI22_X1 _06829_ (.A1(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[29][2] ),
    .A2(net145),
    .B1(net259),
    .B2(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[1][2] ),
    .ZN(_02592_));
 AOI22_X1 _06830_ (.A1(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[23][2] ),
    .A2(net101),
    .B1(net106),
    .B2(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[15][2] ),
    .ZN(_02593_));
 AOI22_X1 _06831_ (.A1(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[2][2] ),
    .A2(net241),
    .B1(net224),
    .B2(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[22][2] ),
    .ZN(_02594_));
 AOI22_X1 _06832_ (.A1(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[16][2] ),
    .A2(net118),
    .B1(net170),
    .B2(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[26][2] ),
    .ZN(_02595_));
 NAND4_X1 _06833_ (.A1(_02592_),
    .A2(_02593_),
    .A3(_02594_),
    .A4(_02595_),
    .ZN(_02596_));
 NOR4_X1 _06834_ (.A1(_02581_),
    .A2(_02586_),
    .A3(_02591_),
    .A4(_02596_),
    .ZN(_02597_));
 OAI21_X1 _06835_ (.A(_01169_),
    .B1(net130),
    .B2(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[0][2] ),
    .ZN(_02598_));
 OAI22_X1 _06836_ (.A1(_02575_),
    .A2(_02576_),
    .B1(_02597_),
    .B2(_02598_),
    .ZN(_02599_));
 NOR4_X1 _06837_ (.A1(_02456_),
    .A2(_02501_),
    .A3(_02546_),
    .A4(_02599_),
    .ZN(_02600_));
 AOI22_X1 _06838_ (.A1(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[26][2] ),
    .A2(net173),
    .B1(net90),
    .B2(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[10][2] ),
    .ZN(_02601_));
 AOI22_X1 _06839_ (.A1(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[3][2] ),
    .A2(net64),
    .B1(net85),
    .B2(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[14][2] ),
    .ZN(_02602_));
 AOI22_X1 _06840_ (.A1(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[8][2] ),
    .A2(net179),
    .B1(net250),
    .B2(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[20][2] ),
    .ZN(_02603_));
 AOI22_X2 _06841_ (.A1(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[27][2] ),
    .A2(net190),
    .B1(net153),
    .B2(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[25][2] ),
    .ZN(_02604_));
 NAND4_X2 _06842_ (.A1(_02601_),
    .A2(_02602_),
    .A3(_02603_),
    .A4(_02604_),
    .ZN(_02605_));
 AOI22_X1 _06843_ (.A1(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[23][2] ),
    .A2(net100),
    .B1(net116),
    .B2(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[16][2] ),
    .ZN(_02606_));
 AOI22_X1 _06844_ (.A1(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[17][2] ),
    .A2(net79),
    .B1(net217),
    .B2(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[9][2] ),
    .ZN(_02607_));
 AOI22_X1 _06845_ (.A1(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[30][2] ),
    .A2(net208),
    .B1(net204),
    .B2(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[13][2] ),
    .ZN(_02608_));
 AOI21_X1 _06846_ (.A(net114),
    .B1(net194),
    .B2(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[19][2] ),
    .ZN(_02609_));
 NAND4_X1 _06847_ (.A1(_02606_),
    .A2(_02607_),
    .A3(_02608_),
    .A4(_02609_),
    .ZN(_02610_));
 AOI22_X1 _06848_ (.A1(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[15][2] ),
    .A2(net107),
    .B1(net93),
    .B2(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[31][2] ),
    .ZN(_02611_));
 AOI22_X1 _06849_ (.A1(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[5][2] ),
    .A2(net131),
    .B1(net82),
    .B2(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[21][2] ),
    .ZN(_02612_));
 AOI22_X1 _06850_ (.A1(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[29][2] ),
    .A2(net142),
    .B1(net255),
    .B2(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[1][2] ),
    .ZN(_02613_));
 AOI22_X1 _06851_ (.A1(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[7][2] ),
    .A2(net68),
    .B1(net233),
    .B2(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[11][2] ),
    .ZN(_02614_));
 NAND4_X1 _06852_ (.A1(_02611_),
    .A2(_02612_),
    .A3(_02613_),
    .A4(_02614_),
    .ZN(_02615_));
 AOI22_X1 _06853_ (.A1(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[24][2] ),
    .A2(net71),
    .B1(net240),
    .B2(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[2][2] ),
    .ZN(_02616_));
 AOI22_X1 _06854_ (.A1(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[4][2] ),
    .A2(net123),
    .B1(net263),
    .B2(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[18][2] ),
    .ZN(_02617_));
 AOI22_X1 _06855_ (.A1(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[12][2] ),
    .A2(net267),
    .B1(net226),
    .B2(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[22][2] ),
    .ZN(_02618_));
 AOI22_X1 _06856_ (.A1(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[28][2] ),
    .A2(net76),
    .B1(net162),
    .B2(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[6][2] ),
    .ZN(_02619_));
 NAND4_X1 _06857_ (.A1(_02616_),
    .A2(_02617_),
    .A3(_02618_),
    .A4(_02619_),
    .ZN(_02620_));
 OR4_X2 _06858_ (.A1(_02605_),
    .A2(_02610_),
    .A3(_02615_),
    .A4(_02620_),
    .ZN(_02621_));
 OAI21_X1 _06859_ (.A(_02621_),
    .B1(net130),
    .B2(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[0][2] ),
    .ZN(_02622_));
 AOI221_X2 _06860_ (.A(_00907_),
    .B1(_02409_),
    .B2(_02600_),
    .C1(_02622_),
    .C2(_01820_),
    .ZN(\rdata_o_n[2] ));
 AOI22_X1 _06861_ (.A1(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[25][3] ),
    .A2(net153),
    .B1(net234),
    .B2(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[11][3] ),
    .ZN(_02623_));
 AOI22_X1 _06862_ (.A1(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[8][3] ),
    .A2(net179),
    .B1(net170),
    .B2(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[26][3] ),
    .ZN(_02624_));
 AOI22_X1 _06863_ (.A1(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[12][3] ),
    .A2(net269),
    .B1(net265),
    .B2(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[18][3] ),
    .ZN(_02625_));
 AOI22_X1 _06864_ (.A1(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[4][3] ),
    .A2(net124),
    .B1(net256),
    .B2(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[1][3] ),
    .ZN(_02626_));
 NAND4_X1 _06865_ (.A1(_02623_),
    .A2(_02624_),
    .A3(_02625_),
    .A4(_02626_),
    .ZN(_02627_));
 AOI22_X1 _06866_ (.A1(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[5][3] ),
    .A2(net132),
    .B1(net226),
    .B2(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[22][3] ),
    .ZN(_02628_));
 AOI22_X1 _06867_ (.A1(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[21][3] ),
    .A2(net82),
    .B1(net219),
    .B2(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[9][3] ),
    .ZN(_02629_));
 AOI22_X1 _06868_ (.A1(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[23][3] ),
    .A2(net101),
    .B1(net251),
    .B2(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[20][3] ),
    .ZN(_02630_));
 AOI21_X1 _06869_ (.A(net113),
    .B1(net190),
    .B2(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[27][3] ),
    .ZN(_02631_));
 NAND4_X1 _06870_ (.A1(_02628_),
    .A2(_02629_),
    .A3(_02630_),
    .A4(_02631_),
    .ZN(_02632_));
 AOI22_X1 _06871_ (.A1(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[31][3] ),
    .A2(net95),
    .B1(net90),
    .B2(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[10][3] ),
    .ZN(_02633_));
 AOI22_X1 _06872_ (.A1(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[15][3] ),
    .A2(net107),
    .B1(net194),
    .B2(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[19][3] ),
    .ZN(_02634_));
 AOI22_X1 _06873_ (.A1(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[28][3] ),
    .A2(net77),
    .B1(net142),
    .B2(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[29][3] ),
    .ZN(_02635_));
 AOI22_X1 _06874_ (.A1(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[17][3] ),
    .A2(net80),
    .B1(net117),
    .B2(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[16][3] ),
    .ZN(_02636_));
 NAND4_X1 _06875_ (.A1(_02633_),
    .A2(_02634_),
    .A3(_02635_),
    .A4(_02636_),
    .ZN(_02637_));
 AOI22_X1 _06876_ (.A1(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[14][3] ),
    .A2(net85),
    .B1(net204),
    .B2(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[13][3] ),
    .ZN(_02638_));
 AOI22_X1 _06877_ (.A1(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[2][3] ),
    .A2(net242),
    .B1(net209),
    .B2(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[30][3] ),
    .ZN(_02639_));
 AOI22_X1 _06878_ (.A1(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[3][3] ),
    .A2(net64),
    .B1(net74),
    .B2(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[24][3] ),
    .ZN(_02640_));
 AOI22_X1 _06879_ (.A1(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[6][3] ),
    .A2(net163),
    .B1(net68),
    .B2(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[7][3] ),
    .ZN(_02641_));
 NAND4_X1 _06880_ (.A1(_02638_),
    .A2(_02639_),
    .A3(_02640_),
    .A4(_02641_),
    .ZN(_02642_));
 NOR4_X1 _06881_ (.A1(_02627_),
    .A2(_02632_),
    .A3(_02637_),
    .A4(_02642_),
    .ZN(_02643_));
 OAI21_X1 _06882_ (.A(_01539_),
    .B1(net130),
    .B2(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[0][3] ),
    .ZN(_02644_));
 AOI22_X1 _06883_ (.A1(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[28][3] ),
    .A2(net77),
    .B1(net193),
    .B2(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[19][3] ),
    .ZN(_02645_));
 AOI22_X1 _06884_ (.A1(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[29][3] ),
    .A2(net144),
    .B1(net132),
    .B2(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[5][3] ),
    .ZN(_02646_));
 AOI22_X1 _06885_ (.A1(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[11][3] ),
    .A2(net236),
    .B1(net212),
    .B2(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[30][3] ),
    .ZN(_02647_));
 AOI22_X1 _06886_ (.A1(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[6][3] ),
    .A2(net163),
    .B1(net68),
    .B2(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[7][3] ),
    .ZN(_02648_));
 NAND4_X1 _06887_ (.A1(_02645_),
    .A2(_02646_),
    .A3(_02647_),
    .A4(_02648_),
    .ZN(_02649_));
 AOI22_X1 _06888_ (.A1(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[21][3] ),
    .A2(net83),
    .B1(net217),
    .B2(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[9][3] ),
    .ZN(_02650_));
 AOI22_X1 _06889_ (.A1(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[17][3] ),
    .A2(net79),
    .B1(net66),
    .B2(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[3][3] ),
    .ZN(_02651_));
 AOI22_X1 _06890_ (.A1(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[22][3] ),
    .A2(net222),
    .B1(net203),
    .B2(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[13][3] ),
    .ZN(_02652_));
 AOI21_X1 _06891_ (.A(net114),
    .B1(net175),
    .B2(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[26][3] ),
    .ZN(_02653_));
 NAND4_X1 _06892_ (.A1(_02650_),
    .A2(_02651_),
    .A3(_02652_),
    .A4(_02653_),
    .ZN(_02654_));
 AOI22_X1 _06893_ (.A1(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[12][3] ),
    .A2(net269),
    .B1(net263),
    .B2(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[18][3] ),
    .ZN(_02655_));
 AOI22_X1 _06894_ (.A1(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[25][3] ),
    .A2(net152),
    .B1(net126),
    .B2(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[4][3] ),
    .ZN(_02656_));
 AOI22_X1 _06895_ (.A1(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[10][3] ),
    .A2(net90),
    .B1(net87),
    .B2(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[14][3] ),
    .ZN(_02657_));
 AOI22_X1 _06896_ (.A1(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[27][3] ),
    .A2(net188),
    .B1(net93),
    .B2(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[31][3] ),
    .ZN(_02658_));
 NAND4_X1 _06897_ (.A1(_02655_),
    .A2(_02656_),
    .A3(_02657_),
    .A4(_02658_),
    .ZN(_02659_));
 AOI22_X1 _06898_ (.A1(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[23][3] ),
    .A2(net104),
    .B1(net260),
    .B2(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[1][3] ),
    .ZN(_02660_));
 AOI22_X1 _06899_ (.A1(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[16][3] ),
    .A2(net117),
    .B1(net242),
    .B2(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[2][3] ),
    .ZN(_02661_));
 AOI22_X1 _06900_ (.A1(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[8][3] ),
    .A2(net180),
    .B1(net245),
    .B2(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[20][3] ),
    .ZN(_02662_));
 AOI22_X1 _06901_ (.A1(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[15][3] ),
    .A2(net108),
    .B1(net71),
    .B2(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[24][3] ),
    .ZN(_02663_));
 NAND4_X1 _06902_ (.A1(_02660_),
    .A2(_02661_),
    .A3(_02662_),
    .A4(_02663_),
    .ZN(_02664_));
 NOR4_X1 _06903_ (.A1(_02649_),
    .A2(_02654_),
    .A3(_02659_),
    .A4(_02664_),
    .ZN(_02665_));
 OAI21_X1 _06904_ (.A(_01700_),
    .B1(net130),
    .B2(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[0][3] ),
    .ZN(_02666_));
 OAI22_X1 _06905_ (.A1(_02643_),
    .A2(_02644_),
    .B1(_02665_),
    .B2(_02666_),
    .ZN(_02667_));
 AOI22_X1 _06906_ (.A1(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[20][3] ),
    .A2(net250),
    .B1(net222),
    .B2(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[22][3] ),
    .ZN(_02668_));
 AOI22_X1 _06907_ (.A1(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[28][3] ),
    .A2(net76),
    .B1(net144),
    .B2(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[29][3] ),
    .ZN(_02669_));
 AOI22_X2 _06908_ (.A1(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[14][3] ),
    .A2(net87),
    .B1(net208),
    .B2(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[30][3] ),
    .ZN(_02670_));
 AOI22_X2 _06909_ (.A1(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[7][3] ),
    .A2(net68),
    .B1(net83),
    .B2(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[21][3] ),
    .ZN(_02671_));
 NAND4_X2 _06910_ (.A1(_02668_),
    .A2(_02669_),
    .A3(_02670_),
    .A4(_02671_),
    .ZN(_02672_));
 AOI22_X1 _06911_ (.A1(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[27][3] ),
    .A2(net188),
    .B1(net204),
    .B2(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[13][3] ),
    .ZN(_02673_));
 AOI22_X1 _06912_ (.A1(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[10][3] ),
    .A2(net90),
    .B1(net254),
    .B2(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[1][3] ),
    .ZN(_02674_));
 AOI22_X1 _06913_ (.A1(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[8][3] ),
    .A2(net180),
    .B1(net267),
    .B2(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[12][3] ),
    .ZN(_02675_));
 AOI21_X1 _06914_ (.A(net114),
    .B1(net236),
    .B2(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[11][3] ),
    .ZN(_02676_));
 NAND4_X1 _06915_ (.A1(_02673_),
    .A2(_02674_),
    .A3(_02675_),
    .A4(_02676_),
    .ZN(_02677_));
 AOI22_X1 _06916_ (.A1(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[3][3] ),
    .A2(net66),
    .B1(net173),
    .B2(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[26][3] ),
    .ZN(_02678_));
 AOI22_X1 _06917_ (.A1(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[16][3] ),
    .A2(net116),
    .B1(net71),
    .B2(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[24][3] ),
    .ZN(_02679_));
 AOI22_X1 _06918_ (.A1(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[25][3] ),
    .A2(net152),
    .B1(net93),
    .B2(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[31][3] ),
    .ZN(_02680_));
 AOI22_X1 _06919_ (.A1(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[2][3] ),
    .A2(net240),
    .B1(net193),
    .B2(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[19][3] ),
    .ZN(_02681_));
 NAND4_X1 _06920_ (.A1(_02678_),
    .A2(_02679_),
    .A3(_02680_),
    .A4(_02681_),
    .ZN(_02682_));
 AOI22_X1 _06921_ (.A1(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[17][3] ),
    .A2(net79),
    .B1(net123),
    .B2(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[4][3] ),
    .ZN(_02683_));
 AOI22_X1 _06922_ (.A1(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[23][3] ),
    .A2(net100),
    .B1(net107),
    .B2(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[15][3] ),
    .ZN(_02684_));
 AOI22_X1 _06923_ (.A1(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[6][3] ),
    .A2(net162),
    .B1(net217),
    .B2(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[9][3] ),
    .ZN(_02685_));
 AOI22_X1 _06924_ (.A1(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[5][3] ),
    .A2(net131),
    .B1(net263),
    .B2(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[18][3] ),
    .ZN(_02686_));
 NAND4_X1 _06925_ (.A1(_02683_),
    .A2(_02684_),
    .A3(_02685_),
    .A4(_02686_),
    .ZN(_02687_));
 NOR4_X1 _06926_ (.A1(_02672_),
    .A2(_02677_),
    .A3(_02682_),
    .A4(_02687_),
    .ZN(_02688_));
 OAI21_X1 _06927_ (.A(_01401_),
    .B1(net130),
    .B2(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[0][3] ),
    .ZN(_02689_));
 OAI21_X1 _06928_ (.A(_01406_),
    .B1(_02688_),
    .B2(_02689_),
    .ZN(_02690_));
 AOI22_X1 _06929_ (.A1(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[31][3] ),
    .A2(net94),
    .B1(net239),
    .B2(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[2][3] ),
    .ZN(_02691_));
 AOI22_X1 _06930_ (.A1(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[18][3] ),
    .A2(_00964_),
    .B1(net200),
    .B2(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[19][3] ),
    .ZN(_02692_));
 AOI22_X1 _06931_ (.A1(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[16][3] ),
    .A2(net121),
    .B1(net88),
    .B2(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[14][3] ),
    .ZN(_02693_));
 AOI22_X2 _06932_ (.A1(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[6][3] ),
    .A2(net159),
    .B1(_00993_),
    .B2(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[11][3] ),
    .ZN(_02694_));
 NAND4_X2 _06933_ (.A1(_02691_),
    .A2(_02692_),
    .A3(_02693_),
    .A4(_02694_),
    .ZN(_02695_));
 AOI22_X1 _06934_ (.A1(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[20][3] ),
    .A2(net246),
    .B1(net216),
    .B2(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[30][3] ),
    .ZN(_02696_));
 AOI22_X1 _06935_ (.A1(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[25][3] ),
    .A2(net151),
    .B1(net141),
    .B2(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[29][3] ),
    .ZN(_02697_));
 AOI22_X1 _06936_ (.A1(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[27][3] ),
    .A2(net186),
    .B1(net129),
    .B2(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[4][3] ),
    .ZN(_02698_));
 AOI21_X1 _06937_ (.A(net115),
    .B1(net89),
    .B2(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[10][3] ),
    .ZN(_02699_));
 NAND4_X2 _06938_ (.A1(_02696_),
    .A2(_02697_),
    .A3(_02698_),
    .A4(_02699_),
    .ZN(_02700_));
 AOI22_X1 _06939_ (.A1(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[23][3] ),
    .A2(_01144_),
    .B1(_01032_),
    .B2(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[28][3] ),
    .ZN(_02701_));
 AOI22_X1 _06940_ (.A1(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[1][3] ),
    .A2(net262),
    .B1(_01007_),
    .B2(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[13][3] ),
    .ZN(_02702_));
 AOI22_X1 _06941_ (.A1(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[24][3] ),
    .A2(_01059_),
    .B1(_00981_),
    .B2(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[21][3] ),
    .ZN(_02703_));
 AOI22_X2 _06942_ (.A1(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[15][3] ),
    .A2(net111),
    .B1(net177),
    .B2(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[8][3] ),
    .ZN(_02704_));
 NAND4_X2 _06943_ (.A1(_02701_),
    .A2(_02702_),
    .A3(_02703_),
    .A4(_02704_),
    .ZN(_02705_));
 AOI22_X1 _06944_ (.A1(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[17][3] ),
    .A2(net81),
    .B1(net221),
    .B2(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[9][3] ),
    .ZN(_02706_));
 AOI22_X1 _06945_ (.A1(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[3][3] ),
    .A2(net63),
    .B1(net167),
    .B2(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[26][3] ),
    .ZN(_02707_));
 AOI22_X1 _06946_ (.A1(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[12][3] ),
    .A2(net274),
    .B1(net227),
    .B2(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[22][3] ),
    .ZN(_02708_));
 AOI22_X1 _06947_ (.A1(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[5][3] ),
    .A2(net135),
    .B1(net70),
    .B2(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[7][3] ),
    .ZN(_02709_));
 NAND4_X2 _06948_ (.A1(_02706_),
    .A2(_02707_),
    .A3(_02708_),
    .A4(_02709_),
    .ZN(_02710_));
 NOR4_X4 _06949_ (.A1(_02695_),
    .A2(_02700_),
    .A3(_02705_),
    .A4(_02710_),
    .ZN(_02711_));
 OAI21_X1 _06950_ (.A(_01662_),
    .B1(net130),
    .B2(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[0][3] ),
    .ZN(_02712_));
 AOI22_X1 _06951_ (.A1(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[3][3] ),
    .A2(net64),
    .B1(net270),
    .B2(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[12][3] ),
    .ZN(_02713_));
 AOI22_X1 _06952_ (.A1(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[27][3] ),
    .A2(net189),
    .B1(net257),
    .B2(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[1][3] ),
    .ZN(_02714_));
 AOI22_X1 _06953_ (.A1(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[15][3] ),
    .A2(net106),
    .B1(net220),
    .B2(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[9][3] ),
    .ZN(_02715_));
 AOI22_X2 _06954_ (.A1(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[29][3] ),
    .A2(net143),
    .B1(net264),
    .B2(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[18][3] ),
    .ZN(_02716_));
 NAND4_X2 _06955_ (.A1(_02713_),
    .A2(_02714_),
    .A3(_02715_),
    .A4(_02716_),
    .ZN(_02717_));
 AOI22_X1 _06956_ (.A1(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[26][3] ),
    .A2(net168),
    .B1(net136),
    .B2(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[5][3] ),
    .ZN(_02718_));
 AOI22_X1 _06957_ (.A1(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[8][3] ),
    .A2(net183),
    .B1(net125),
    .B2(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[4][3] ),
    .ZN(_02719_));
 AOI22_X1 _06958_ (.A1(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[10][3] ),
    .A2(net91),
    .B1(net197),
    .B2(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[19][3] ),
    .ZN(_02720_));
 AOI21_X1 _06959_ (.A(_01119_),
    .B1(net96),
    .B2(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[31][3] ),
    .ZN(_02721_));
 NAND4_X2 _06960_ (.A1(_02718_),
    .A2(_02719_),
    .A3(_02720_),
    .A4(_02721_),
    .ZN(_02722_));
 AOI22_X1 _06961_ (.A1(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[16][3] ),
    .A2(net118),
    .B1(net67),
    .B2(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[7][3] ),
    .ZN(_02723_));
 AOI22_X1 _06962_ (.A1(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[17][3] ),
    .A2(net80),
    .B1(net82),
    .B2(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[21][3] ),
    .ZN(_02724_));
 AOI22_X1 _06963_ (.A1(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[2][3] ),
    .A2(net243),
    .B1(net225),
    .B2(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[22][3] ),
    .ZN(_02725_));
 AOI22_X1 _06964_ (.A1(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[28][3] ),
    .A2(net75),
    .B1(net161),
    .B2(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[6][3] ),
    .ZN(_02726_));
 NAND4_X2 _06965_ (.A1(_02723_),
    .A2(_02724_),
    .A3(_02725_),
    .A4(_02726_),
    .ZN(_02727_));
 AOI22_X1 _06966_ (.A1(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[23][3] ),
    .A2(net103),
    .B1(net72),
    .B2(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[24][3] ),
    .ZN(_02728_));
 AOI22_X1 _06967_ (.A1(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[20][3] ),
    .A2(net247),
    .B1(net210),
    .B2(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[30][3] ),
    .ZN(_02729_));
 AOI22_X1 _06968_ (.A1(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[11][3] ),
    .A2(net232),
    .B1(net206),
    .B2(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[13][3] ),
    .ZN(_02730_));
 AOI22_X2 _06969_ (.A1(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[25][3] ),
    .A2(net154),
    .B1(net86),
    .B2(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[14][3] ),
    .ZN(_02731_));
 NAND4_X2 _06970_ (.A1(_02728_),
    .A2(_02729_),
    .A3(_02730_),
    .A4(_02731_),
    .ZN(_02732_));
 NOR4_X4 _06971_ (.A1(_02717_),
    .A2(_02722_),
    .A3(_02727_),
    .A4(_02732_),
    .ZN(_02733_));
 OAI21_X1 _06972_ (.A(_01164_),
    .B1(net130),
    .B2(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[0][3] ),
    .ZN(_02734_));
 OAI22_X1 _06973_ (.A1(_02711_),
    .A2(_02712_),
    .B1(_02733_),
    .B2(_02734_),
    .ZN(_02735_));
 AOI22_X1 _06974_ (.A1(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[8][3] ),
    .A2(net176),
    .B1(_01007_),
    .B2(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[13][3] ),
    .ZN(_02736_));
 AOI22_X1 _06975_ (.A1(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[5][3] ),
    .A2(net135),
    .B1(net70),
    .B2(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[7][3] ),
    .ZN(_02737_));
 AOI22_X1 _06976_ (.A1(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[15][3] ),
    .A2(net111),
    .B1(net221),
    .B2(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[9][3] ),
    .ZN(_02738_));
 AOI22_X2 _06977_ (.A1(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[3][3] ),
    .A2(net63),
    .B1(net159),
    .B2(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[6][3] ),
    .ZN(_02739_));
 NAND4_X2 _06978_ (.A1(_02736_),
    .A2(_02737_),
    .A3(_02738_),
    .A4(_02739_),
    .ZN(_02740_));
 AOI22_X1 _06979_ (.A1(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[26][3] ),
    .A2(net167),
    .B1(net89),
    .B2(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[10][3] ),
    .ZN(_02741_));
 AOI22_X1 _06980_ (.A1(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[27][3] ),
    .A2(net186),
    .B1(net121),
    .B2(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[16][3] ),
    .ZN(_02742_));
 AOI22_X1 _06981_ (.A1(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[23][3] ),
    .A2(_01144_),
    .B1(net151),
    .B2(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[25][3] ),
    .ZN(_02743_));
 AOI21_X1 _06982_ (.A(net115),
    .B1(_00996_),
    .B2(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[22][3] ),
    .ZN(_02744_));
 NAND4_X2 _06983_ (.A1(_02741_),
    .A2(_02742_),
    .A3(_02743_),
    .A4(_02744_),
    .ZN(_02745_));
 AOI22_X1 _06984_ (.A1(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[29][3] ),
    .A2(_01050_),
    .B1(net231),
    .B2(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[11][3] ),
    .ZN(_02746_));
 AOI22_X1 _06985_ (.A1(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[28][3] ),
    .A2(_01032_),
    .B1(net200),
    .B2(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[19][3] ),
    .ZN(_02747_));
 AOI22_X1 _06986_ (.A1(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[17][3] ),
    .A2(net81),
    .B1(net244),
    .B2(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[20][3] ),
    .ZN(_02748_));
 AOI22_X2 _06987_ (.A1(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[21][3] ),
    .A2(_00981_),
    .B1(net215),
    .B2(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[30][3] ),
    .ZN(_02749_));
 NAND4_X2 _06988_ (.A1(_02746_),
    .A2(_02747_),
    .A3(_02748_),
    .A4(_02749_),
    .ZN(_02750_));
 AOI22_X1 _06989_ (.A1(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[24][3] ),
    .A2(_01059_),
    .B1(net88),
    .B2(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[14][3] ),
    .ZN(_02751_));
 AOI22_X1 _06990_ (.A1(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[12][3] ),
    .A2(net274),
    .B1(net262),
    .B2(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[1][3] ),
    .ZN(_02752_));
 AOI22_X1 _06991_ (.A1(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[31][3] ),
    .A2(_01149_),
    .B1(_00964_),
    .B2(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[18][3] ),
    .ZN(_02753_));
 AOI22_X2 _06992_ (.A1(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[4][3] ),
    .A2(net129),
    .B1(_00989_),
    .B2(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[2][3] ),
    .ZN(_02754_));
 NAND4_X2 _06993_ (.A1(_02751_),
    .A2(_02752_),
    .A3(_02753_),
    .A4(_02754_),
    .ZN(_02755_));
 NOR4_X4 _06994_ (.A1(_02740_),
    .A2(_02745_),
    .A3(_02750_),
    .A4(_02755_),
    .ZN(_02756_));
 OAI21_X1 _06995_ (.A(_01502_),
    .B1(net130),
    .B2(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[0][3] ),
    .ZN(_02757_));
 AOI22_X1 _06996_ (.A1(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[4][3] ),
    .A2(net125),
    .B1(net235),
    .B2(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[11][3] ),
    .ZN(_02758_));
 AOI22_X1 _06997_ (.A1(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[8][3] ),
    .A2(_01034_),
    .B1(net68),
    .B2(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[7][3] ),
    .ZN(_02759_));
 AOI22_X1 _06998_ (.A1(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[26][3] ),
    .A2(_01038_),
    .B1(net205),
    .B2(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[13][3] ),
    .ZN(_02760_));
 AOI22_X1 _06999_ (.A1(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[23][3] ),
    .A2(net105),
    .B1(net241),
    .B2(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[2][3] ),
    .ZN(_02761_));
 NAND4_X1 _07000_ (.A1(_02758_),
    .A2(_02759_),
    .A3(_02760_),
    .A4(_02761_),
    .ZN(_02762_));
 AOI22_X1 _07001_ (.A1(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[3][3] ),
    .A2(net65),
    .B1(net86),
    .B2(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[14][3] ),
    .ZN(_02763_));
 AOI22_X1 _07002_ (.A1(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[31][3] ),
    .A2(net96),
    .B1(net220),
    .B2(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[9][3] ),
    .ZN(_02764_));
 AOI22_X1 _07003_ (.A1(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[10][3] ),
    .A2(net91),
    .B1(net225),
    .B2(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[22][3] ),
    .ZN(_02765_));
 AOI21_X1 _07004_ (.A(net113),
    .B1(net155),
    .B2(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[25][3] ),
    .ZN(_02766_));
 NAND4_X1 _07005_ (.A1(_02763_),
    .A2(_02764_),
    .A3(_02765_),
    .A4(_02766_),
    .ZN(_02767_));
 AOI22_X1 _07006_ (.A1(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[5][3] ),
    .A2(net138),
    .B1(_01009_),
    .B2(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[19][3] ),
    .ZN(_02768_));
 AOI22_X1 _07007_ (.A1(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[21][3] ),
    .A2(net83),
    .B1(net211),
    .B2(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[30][3] ),
    .ZN(_02769_));
 AOI22_X1 _07008_ (.A1(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[16][3] ),
    .A2(_01097_),
    .B1(net249),
    .B2(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[20][3] ),
    .ZN(_02770_));
 AOI22_X1 _07009_ (.A1(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[29][3] ),
    .A2(net145),
    .B1(net72),
    .B2(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[24][3] ),
    .ZN(_02771_));
 NAND4_X1 _07010_ (.A1(_02768_),
    .A2(_02769_),
    .A3(_02770_),
    .A4(_02771_),
    .ZN(_02772_));
 AOI22_X1 _07011_ (.A1(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[27][3] ),
    .A2(net192),
    .B1(net77),
    .B2(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[28][3] ),
    .ZN(_02773_));
 AOI22_X1 _07012_ (.A1(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[6][3] ),
    .A2(net164),
    .B1(net260),
    .B2(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[1][3] ),
    .ZN(_02774_));
 AOI22_X1 _07013_ (.A1(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[17][3] ),
    .A2(net78),
    .B1(net108),
    .B2(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[15][3] ),
    .ZN(_02775_));
 AOI22_X1 _07014_ (.A1(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[12][3] ),
    .A2(net271),
    .B1(net265),
    .B2(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[18][3] ),
    .ZN(_02776_));
 NAND4_X1 _07015_ (.A1(_02773_),
    .A2(_02774_),
    .A3(_02775_),
    .A4(_02776_),
    .ZN(_02777_));
 NOR4_X1 _07016_ (.A1(_02762_),
    .A2(_02767_),
    .A3(_02772_),
    .A4(_02777_),
    .ZN(_02778_));
 OAI21_X1 _07017_ (.A(_01764_),
    .B1(net130),
    .B2(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[0][3] ),
    .ZN(_02779_));
 OAI22_X2 _07018_ (.A1(_02756_),
    .A2(_02757_),
    .B1(_02778_),
    .B2(_02779_),
    .ZN(_02780_));
 NOR4_X1 _07019_ (.A1(_02667_),
    .A2(_02690_),
    .A3(_02735_),
    .A4(_02780_),
    .ZN(_02781_));
 AOI22_X1 _07020_ (.A1(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[25][3] ),
    .A2(net147),
    .B1(net218),
    .B2(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[9][3] ),
    .ZN(_02782_));
 AOI22_X1 _07021_ (.A1(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[4][3] ),
    .A2(net127),
    .B1(net203),
    .B2(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[13][3] ),
    .ZN(_02783_));
 AOI22_X1 _07022_ (.A1(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[15][3] ),
    .A2(net110),
    .B1(net202),
    .B2(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[19][3] ),
    .ZN(_02784_));
 AOI22_X1 _07023_ (.A1(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[18][3] ),
    .A2(_00964_),
    .B1(net230),
    .B2(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[11][3] ),
    .ZN(_02785_));
 NAND4_X1 _07024_ (.A1(_02782_),
    .A2(_02783_),
    .A3(_02784_),
    .A4(_02785_),
    .ZN(_02786_));
 AOI22_X1 _07025_ (.A1(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[29][3] ),
    .A2(net141),
    .B1(net94),
    .B2(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[31][3] ),
    .ZN(_02787_));
 AOI22_X1 _07026_ (.A1(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[5][3] ),
    .A2(net133),
    .B1(_01059_),
    .B2(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[24][3] ),
    .ZN(_02788_));
 MUX2_X1 _07027_ (.A(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[12][3] ),
    .B(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[14][3] ),
    .S(net8),
    .Z(_02789_));
 AOI221_X1 _07028_ (.A(net115),
    .B1(net92),
    .B2(_02789_),
    .C1(net214),
    .C2(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[30][3] ),
    .ZN(_02790_));
 NAND3_X1 _07029_ (.A1(_02787_),
    .A2(_02788_),
    .A3(_02790_),
    .ZN(_02791_));
 AOI22_X1 _07030_ (.A1(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[3][3] ),
    .A2(net63),
    .B1(net177),
    .B2(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[8][3] ),
    .ZN(_02792_));
 AOI22_X1 _07031_ (.A1(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[23][3] ),
    .A2(net97),
    .B1(net122),
    .B2(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[16][3] ),
    .ZN(_02793_));
 AOI22_X1 _07032_ (.A1(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[20][3] ),
    .A2(net246),
    .B1(net227),
    .B2(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[22][3] ),
    .ZN(_02794_));
 AOI22_X2 _07033_ (.A1(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[6][3] ),
    .A2(net159),
    .B1(net239),
    .B2(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[2][3] ),
    .ZN(_02795_));
 NAND4_X2 _07034_ (.A1(_02792_),
    .A2(_02793_),
    .A3(_02794_),
    .A4(_02795_),
    .ZN(_02796_));
 AOI22_X1 _07035_ (.A1(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[10][3] ),
    .A2(_00956_),
    .B1(net261),
    .B2(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[1][3] ),
    .ZN(_02797_));
 AOI22_X1 _07036_ (.A1(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[17][3] ),
    .A2(net81),
    .B1(net69),
    .B2(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[7][3] ),
    .ZN(_02798_));
 AOI22_X1 _07037_ (.A1(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[28][3] ),
    .A2(net76),
    .B1(net166),
    .B2(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[26][3] ),
    .ZN(_02799_));
 AOI22_X1 _07038_ (.A1(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[27][3] ),
    .A2(net187),
    .B1(_00981_),
    .B2(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[21][3] ),
    .ZN(_02800_));
 NAND4_X1 _07039_ (.A1(_02797_),
    .A2(_02798_),
    .A3(_02799_),
    .A4(_02800_),
    .ZN(_02801_));
 NOR4_X2 _07040_ (.A1(_02786_),
    .A2(_02791_),
    .A3(_02796_),
    .A4(_02801_),
    .ZN(_02802_));
 OAI21_X2 _07041_ (.A(_01623_),
    .B1(net130),
    .B2(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[0][3] ),
    .ZN(_02803_));
 INV_X1 _07042_ (.A(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[27][3] ),
    .ZN(_02804_));
 INV_X1 _07043_ (.A(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[22][3] ),
    .ZN(_02805_));
 OAI22_X1 _07044_ (.A1(_02804_),
    .A2(_02555_),
    .B1(_01216_),
    .B2(_02805_),
    .ZN(_02806_));
 AOI221_X2 _07045_ (.A(_02806_),
    .B1(net263),
    .B2(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[18][3] ),
    .C1(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[28][3] ),
    .C2(net76),
    .ZN(_02807_));
 INV_X1 _07046_ (.A(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[29][3] ),
    .ZN(_02808_));
 INV_X1 _07047_ (.A(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[9][3] ),
    .ZN(_02809_));
 OAI22_X1 _07048_ (.A1(_02808_),
    .A2(_01425_),
    .B1(_01420_),
    .B2(_02809_),
    .ZN(_02810_));
 AOI221_X2 _07049_ (.A(_02810_),
    .B1(net126),
    .B2(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[4][3] ),
    .C1(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[17][3] ),
    .C2(net79),
    .ZN(_02811_));
 INV_X1 _07050_ (.A(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[3][3] ),
    .ZN(_02812_));
 INV_X1 _07051_ (.A(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[24][3] ),
    .ZN(_02813_));
 OAI33_X1 _07052_ (.A1(_02812_),
    .A2(_01015_),
    .A3(_00952_),
    .B1(_00954_),
    .B2(_00979_),
    .B3(_02813_),
    .ZN(_02814_));
 AOI221_X2 _07053_ (.A(_02814_),
    .B1(_00956_),
    .B2(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[10][3] ),
    .C1(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[31][3] ),
    .C2(net93),
    .ZN(_02815_));
 MUX2_X1 _07054_ (.A(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[12][3] ),
    .B(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[14][3] ),
    .S(net8),
    .Z(_02816_));
 AOI221_X2 _07055_ (.A(net114),
    .B1(net92),
    .B2(_02816_),
    .C1(net174),
    .C2(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[26][3] ),
    .ZN(_02817_));
 NAND4_X2 _07056_ (.A1(_02807_),
    .A2(_02811_),
    .A3(_02815_),
    .A4(_02817_),
    .ZN(_02818_));
 AOI22_X1 _07057_ (.A1(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[11][3] ),
    .A2(net229),
    .B1(net203),
    .B2(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[13][3] ),
    .ZN(_02819_));
 AOI22_X1 _07058_ (.A1(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[25][3] ),
    .A2(net148),
    .B1(net196),
    .B2(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[19][3] ),
    .ZN(_02820_));
 AOI22_X1 _07059_ (.A1(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[8][3] ),
    .A2(net178),
    .B1(net238),
    .B2(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[2][3] ),
    .ZN(_02821_));
 AOI22_X1 _07060_ (.A1(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[15][3] ),
    .A2(net110),
    .B1(net134),
    .B2(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[5][3] ),
    .ZN(_02822_));
 NAND4_X1 _07061_ (.A1(_02819_),
    .A2(_02820_),
    .A3(_02821_),
    .A4(_02822_),
    .ZN(_02823_));
 AOI22_X1 _07062_ (.A1(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[1][3] ),
    .A2(net254),
    .B1(net213),
    .B2(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[30][3] ),
    .ZN(_02824_));
 AOI22_X1 _07063_ (.A1(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[16][3] ),
    .A2(net120),
    .B1(net83),
    .B2(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[21][3] ),
    .ZN(_02825_));
 AOI22_X1 _07064_ (.A1(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[6][3] ),
    .A2(net158),
    .B1(net69),
    .B2(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[7][3] ),
    .ZN(_02826_));
 AOI22_X1 _07065_ (.A1(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[23][3] ),
    .A2(net102),
    .B1(net245),
    .B2(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[20][3] ),
    .ZN(_02827_));
 NAND4_X1 _07066_ (.A1(_02824_),
    .A2(_02825_),
    .A3(_02826_),
    .A4(_02827_),
    .ZN(_02828_));
 NOR3_X2 _07067_ (.A1(_02818_),
    .A2(_02823_),
    .A3(_02828_),
    .ZN(_02829_));
 OAI21_X1 _07068_ (.A(_01295_),
    .B1(net130),
    .B2(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[0][3] ),
    .ZN(_02830_));
 OAI22_X4 _07069_ (.A1(_02802_),
    .A2(_02803_),
    .B1(_02829_),
    .B2(_02830_),
    .ZN(_02831_));
 AOI22_X1 _07070_ (.A1(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[29][3] ),
    .A2(net140),
    .B1(net136),
    .B2(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[5][3] ),
    .ZN(_02832_));
 AOI22_X1 _07071_ (.A1(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[15][3] ),
    .A2(net109),
    .B1(net72),
    .B2(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[24][3] ),
    .ZN(_02833_));
 AOI22_X1 _07072_ (.A1(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[7][3] ),
    .A2(net67),
    .B1(net243),
    .B2(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[2][3] ),
    .ZN(_02834_));
 AOI22_X1 _07073_ (.A1(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[23][3] ),
    .A2(net98),
    .B1(net266),
    .B2(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[12][3] ),
    .ZN(_02835_));
 NAND4_X1 _07074_ (.A1(_02832_),
    .A2(_02833_),
    .A3(_02834_),
    .A4(_02835_),
    .ZN(_02836_));
 AOI22_X1 _07075_ (.A1(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[8][3] ),
    .A2(net182),
    .B1(net248),
    .B2(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[20][3] ),
    .ZN(_02837_));
 AOI22_X1 _07076_ (.A1(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[27][3] ),
    .A2(net191),
    .B1(net91),
    .B2(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[10][3] ),
    .ZN(_02838_));
 AOI22_X1 _07077_ (.A1(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[16][3] ),
    .A2(net119),
    .B1(_01149_),
    .B2(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[31][3] ),
    .ZN(_02839_));
 AOI21_X1 _07078_ (.A(_01119_),
    .B1(net207),
    .B2(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[30][3] ),
    .ZN(_02840_));
 NAND4_X2 _07079_ (.A1(_02837_),
    .A2(_02838_),
    .A3(_02839_),
    .A4(_02840_),
    .ZN(_02841_));
 AOI22_X1 _07080_ (.A1(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[26][3] ),
    .A2(net168),
    .B1(net223),
    .B2(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[22][3] ),
    .ZN(_02842_));
 AOI22_X1 _07081_ (.A1(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[17][3] ),
    .A2(net78),
    .B1(net220),
    .B2(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[9][3] ),
    .ZN(_02843_));
 AOI22_X1 _07082_ (.A1(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[21][3] ),
    .A2(net84),
    .B1(net206),
    .B2(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[13][3] ),
    .ZN(_02844_));
 AOI22_X2 _07083_ (.A1(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[3][3] ),
    .A2(net65),
    .B1(net75),
    .B2(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[28][3] ),
    .ZN(_02845_));
 NAND4_X2 _07084_ (.A1(_02842_),
    .A2(_02843_),
    .A3(_02844_),
    .A4(_02845_),
    .ZN(_02846_));
 AOI22_X1 _07085_ (.A1(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[14][3] ),
    .A2(net86),
    .B1(net258),
    .B2(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[1][3] ),
    .ZN(_02847_));
 AOI22_X1 _07086_ (.A1(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[25][3] ),
    .A2(net149),
    .B1(net198),
    .B2(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[19][3] ),
    .ZN(_02848_));
 AOI22_X1 _07087_ (.A1(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[6][3] ),
    .A2(net160),
    .B1(net264),
    .B2(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[18][3] ),
    .ZN(_02849_));
 AOI22_X2 _07088_ (.A1(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[4][3] ),
    .A2(net128),
    .B1(net232),
    .B2(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[11][3] ),
    .ZN(_02850_));
 NAND4_X2 _07089_ (.A1(_02847_),
    .A2(_02848_),
    .A3(_02849_),
    .A4(_02850_),
    .ZN(_02851_));
 NOR4_X2 _07090_ (.A1(_02836_),
    .A2(_02841_),
    .A3(_02846_),
    .A4(_02851_),
    .ZN(_02852_));
 OAI21_X1 _07091_ (.A(_00923_),
    .B1(_01064_),
    .B2(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[0][3] ),
    .ZN(_02853_));
 AOI22_X1 _07092_ (.A1(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[8][3] ),
    .A2(net176),
    .B1(net172),
    .B2(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[26][3] ),
    .ZN(_02854_));
 AOI22_X1 _07093_ (.A1(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[5][3] ),
    .A2(net135),
    .B1(net200),
    .B2(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[19][3] ),
    .ZN(_02855_));
 AND2_X1 _07094_ (.A1(_02854_),
    .A2(_02855_),
    .ZN(_02856_));
 INV_X1 _07095_ (.A(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[15][3] ),
    .ZN(_02857_));
 INV_X1 _07096_ (.A(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[9][3] ),
    .ZN(_02858_));
 OAI22_X1 _07097_ (.A1(_02857_),
    .A2(_01029_),
    .B1(_01420_),
    .B2(_02858_),
    .ZN(_02859_));
 AOI221_X1 _07098_ (.A(_02859_),
    .B1(net63),
    .B2(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[3][3] ),
    .C1(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[16][3] ),
    .C2(net121),
    .ZN(_02860_));
 AOI222_X2 _07099_ (.A1(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[23][3] ),
    .A2(net99),
    .B1(net274),
    .B2(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[12][3] ),
    .C1(net146),
    .C2(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[29][3] ),
    .ZN(_02861_));
 INV_X1 _07100_ (.A(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[17][3] ),
    .ZN(_02862_));
 INV_X1 _07101_ (.A(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[2][3] ),
    .ZN(_02863_));
 OAI33_X1 _07102_ (.A1(_02862_),
    .A2(_01015_),
    .A3(_00979_),
    .B1(_00952_),
    .B2(_00962_),
    .B3(_02863_),
    .ZN(_02864_));
 AOI221_X1 _07103_ (.A(_02864_),
    .B1(net244),
    .B2(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[20][3] ),
    .C1(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[28][3] ),
    .C2(_01032_),
    .ZN(_02865_));
 NAND4_X1 _07104_ (.A1(_02856_),
    .A2(_02860_),
    .A3(_02861_),
    .A4(_02865_),
    .ZN(_02866_));
 AOI221_X1 _07105_ (.A(net115),
    .B1(net89),
    .B2(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[10][3] ),
    .C1(net228),
    .C2(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[22][3] ),
    .ZN(_02867_));
 AOI22_X1 _07106_ (.A1(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[4][3] ),
    .A2(net128),
    .B1(_00971_),
    .B2(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[14][3] ),
    .ZN(_02868_));
 AOI22_X1 _07107_ (.A1(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[6][3] ),
    .A2(net156),
    .B1(net264),
    .B2(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[18][3] ),
    .ZN(_02869_));
 AOI22_X1 _07108_ (.A1(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[24][3] ),
    .A2(net73),
    .B1(_00981_),
    .B2(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[21][3] ),
    .ZN(_02870_));
 NAND4_X1 _07109_ (.A1(_02867_),
    .A2(_02868_),
    .A3(_02869_),
    .A4(_02870_),
    .ZN(_02871_));
 AOI22_X1 _07110_ (.A1(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[25][3] ),
    .A2(net150),
    .B1(net215),
    .B2(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[30][3] ),
    .ZN(_02872_));
 AOI22_X1 _07111_ (.A1(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[7][3] ),
    .A2(net70),
    .B1(net206),
    .B2(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[13][3] ),
    .ZN(_02873_));
 AOI22_X1 _07112_ (.A1(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[27][3] ),
    .A2(_01021_),
    .B1(net237),
    .B2(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[11][3] ),
    .ZN(_02874_));
 AOI22_X2 _07113_ (.A1(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[31][3] ),
    .A2(_01149_),
    .B1(net253),
    .B2(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[1][3] ),
    .ZN(_02875_));
 NAND4_X2 _07114_ (.A1(_02872_),
    .A2(_02873_),
    .A3(_02874_),
    .A4(_02875_),
    .ZN(_02876_));
 NOR3_X2 _07115_ (.A1(_02866_),
    .A2(_02871_),
    .A3(_02876_),
    .ZN(_02877_));
 OAI21_X1 _07116_ (.A(_01731_),
    .B1(_01064_),
    .B2(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[0][3] ),
    .ZN(_02878_));
 OAI22_X2 _07117_ (.A1(_02852_),
    .A2(_02853_),
    .B1(_02877_),
    .B2(_02878_),
    .ZN(_02879_));
 AOI22_X1 _07118_ (.A1(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[16][3] ),
    .A2(net119),
    .B1(_01032_),
    .B2(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[28][3] ),
    .ZN(_02880_));
 AOI22_X1 _07119_ (.A1(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[3][3] ),
    .A2(net65),
    .B1(net252),
    .B2(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[20][3] ),
    .ZN(_02881_));
 AOI22_X1 _07120_ (.A1(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[5][3] ),
    .A2(net139),
    .B1(net237),
    .B2(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[11][3] ),
    .ZN(_02882_));
 AOI22_X1 _07121_ (.A1(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[27][3] ),
    .A2(net192),
    .B1(net73),
    .B2(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[24][3] ),
    .ZN(_02883_));
 NAND4_X1 _07122_ (.A1(_02880_),
    .A2(_02881_),
    .A3(_02882_),
    .A4(_02883_),
    .ZN(_02884_));
 AOI22_X1 _07123_ (.A1(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[6][3] ),
    .A2(net160),
    .B1(net87),
    .B2(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[14][3] ),
    .ZN(_02885_));
 AOI22_X1 _07124_ (.A1(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[23][3] ),
    .A2(net99),
    .B1(net109),
    .B2(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[15][3] ),
    .ZN(_02886_));
 AOI22_X1 _07125_ (.A1(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[17][3] ),
    .A2(net78),
    .B1(net225),
    .B2(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[22][3] ),
    .ZN(_02887_));
 AOI21_X1 _07126_ (.A(_01119_),
    .B1(_01149_),
    .B2(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[31][3] ),
    .ZN(_02888_));
 NAND4_X2 _07127_ (.A1(_02885_),
    .A2(_02886_),
    .A3(_02887_),
    .A4(_02888_),
    .ZN(_02889_));
 AOI22_X1 _07128_ (.A1(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[8][3] ),
    .A2(net183),
    .B1(net264),
    .B2(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[18][3] ),
    .ZN(_02890_));
 AOI22_X1 _07129_ (.A1(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[12][3] ),
    .A2(net272),
    .B1(net89),
    .B2(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[10][3] ),
    .ZN(_02891_));
 AOI22_X1 _07130_ (.A1(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[26][3] ),
    .A2(net171),
    .B1(net243),
    .B2(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[2][3] ),
    .ZN(_02892_));
 AOI22_X1 _07131_ (.A1(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[1][3] ),
    .A2(net253),
    .B1(net198),
    .B2(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[19][3] ),
    .ZN(_02893_));
 NAND4_X1 _07132_ (.A1(_02890_),
    .A2(_02891_),
    .A3(_02892_),
    .A4(_02893_),
    .ZN(_02894_));
 AOI22_X1 _07133_ (.A1(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[30][3] ),
    .A2(net211),
    .B1(net206),
    .B2(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[13][3] ),
    .ZN(_02895_));
 AOI22_X1 _07134_ (.A1(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[21][3] ),
    .A2(net84),
    .B1(_00999_),
    .B2(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[9][3] ),
    .ZN(_02896_));
 AOI22_X1 _07135_ (.A1(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[7][3] ),
    .A2(net70),
    .B1(net128),
    .B2(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[4][3] ),
    .ZN(_02897_));
 AOI22_X2 _07136_ (.A1(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[25][3] ),
    .A2(net150),
    .B1(net146),
    .B2(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[29][3] ),
    .ZN(_02898_));
 NAND4_X2 _07137_ (.A1(_02895_),
    .A2(_02896_),
    .A3(_02897_),
    .A4(_02898_),
    .ZN(_02899_));
 NOR4_X2 _07138_ (.A1(_02884_),
    .A2(_02889_),
    .A3(_02894_),
    .A4(_02899_),
    .ZN(_02900_));
 OAI21_X1 _07139_ (.A(_01408_),
    .B1(net130),
    .B2(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[0][3] ),
    .ZN(_02901_));
 AOI22_X1 _07140_ (.A1(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[3][3] ),
    .A2(_01102_),
    .B1(net76),
    .B2(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[28][3] ),
    .ZN(_02902_));
 AOI22_X1 _07141_ (.A1(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[10][3] ),
    .A2(_00956_),
    .B1(net199),
    .B2(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[19][3] ),
    .ZN(_02903_));
 AOI22_X1 _07142_ (.A1(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[6][3] ),
    .A2(net157),
    .B1(net69),
    .B2(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[7][3] ),
    .ZN(_02904_));
 AOI22_X2 _07143_ (.A1(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[12][3] ),
    .A2(net273),
    .B1(_00964_),
    .B2(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[18][3] ),
    .ZN(_02905_));
 NAND4_X2 _07144_ (.A1(_02902_),
    .A2(_02903_),
    .A3(_02904_),
    .A4(_02905_),
    .ZN(_02906_));
 AOI22_X1 _07145_ (.A1(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[27][3] ),
    .A2(net187),
    .B1(net122),
    .B2(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[16][3] ),
    .ZN(_02907_));
 AOI22_X1 _07146_ (.A1(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[29][3] ),
    .A2(net141),
    .B1(net214),
    .B2(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[30][3] ),
    .ZN(_02908_));
 MUX2_X1 _07147_ (.A(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[24][3] ),
    .B(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[26][3] ),
    .S(net8),
    .Z(_02909_));
 AOI22_X1 _07148_ (.A1(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[8][3] ),
    .A2(_00939_),
    .B1(_02909_),
    .B2(net1),
    .ZN(_02910_));
 INV_X1 _07149_ (.A(_02910_),
    .ZN(_02911_));
 NOR3_X4 _07150_ (.A1(net7),
    .A2(_00944_),
    .A3(net9),
    .ZN(_02912_));
 AOI221_X2 _07151_ (.A(net115),
    .B1(net94),
    .B2(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[31][3] ),
    .C1(_02911_),
    .C2(_02912_),
    .ZN(_02913_));
 NAND3_X2 _07152_ (.A1(_02907_),
    .A2(_02908_),
    .A3(_02913_),
    .ZN(_02914_));
 AOI22_X1 _07153_ (.A1(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[2][3] ),
    .A2(net238),
    .B1(net229),
    .B2(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[11][3] ),
    .ZN(_02915_));
 AOI22_X1 _07154_ (.A1(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[23][3] ),
    .A2(net97),
    .B1(net88),
    .B2(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[14][3] ),
    .ZN(_02916_));
 AOI22_X1 _07155_ (.A1(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[5][3] ),
    .A2(net133),
    .B1(net203),
    .B2(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[13][3] ),
    .ZN(_02917_));
 AOI22_X2 _07156_ (.A1(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[15][3] ),
    .A2(net110),
    .B1(net127),
    .B2(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[4][3] ),
    .ZN(_02918_));
 NAND4_X2 _07157_ (.A1(_02915_),
    .A2(_02916_),
    .A3(_02917_),
    .A4(_02918_),
    .ZN(_02919_));
 AOI222_X2 _07158_ (.A1(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[17][3] ),
    .A2(net81),
    .B1(_00981_),
    .B2(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[21][3] ),
    .C1(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[22][3] ),
    .C2(net227),
    .ZN(_02920_));
 AOI22_X1 _07159_ (.A1(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[25][3] ),
    .A2(net147),
    .B1(net246),
    .B2(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[20][3] ),
    .ZN(_02921_));
 AOI22_X1 _07160_ (.A1(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[1][3] ),
    .A2(net261),
    .B1(net218),
    .B2(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[9][3] ),
    .ZN(_02922_));
 NAND3_X1 _07161_ (.A1(_02920_),
    .A2(_02921_),
    .A3(_02922_),
    .ZN(_02923_));
 NOR4_X4 _07162_ (.A1(_02906_),
    .A2(_02914_),
    .A3(_02919_),
    .A4(_02923_),
    .ZN(_02924_));
 OAI21_X1 _07163_ (.A(_01583_),
    .B1(net130),
    .B2(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[0][3] ),
    .ZN(_02925_));
 OAI22_X2 _07164_ (.A1(_02900_),
    .A2(_02901_),
    .B1(_02924_),
    .B2(_02925_),
    .ZN(_02926_));
 AOI22_X1 _07165_ (.A1(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[25][3] ),
    .A2(net154),
    .B1(net225),
    .B2(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[22][3] ),
    .ZN(_02927_));
 AOI22_X1 _07166_ (.A1(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[3][3] ),
    .A2(net64),
    .B1(net257),
    .B2(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[1][3] ),
    .ZN(_02928_));
 AOI22_X1 _07167_ (.A1(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[24][3] ),
    .A2(net72),
    .B1(net85),
    .B2(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[14][3] ),
    .ZN(_02929_));
 AOI22_X2 _07168_ (.A1(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[27][3] ),
    .A2(net189),
    .B1(net197),
    .B2(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[19][3] ),
    .ZN(_02930_));
 NAND4_X2 _07169_ (.A1(_02927_),
    .A2(_02928_),
    .A3(_02929_),
    .A4(_02930_),
    .ZN(_02931_));
 AOI22_X1 _07170_ (.A1(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[6][3] ),
    .A2(net161),
    .B1(net219),
    .B2(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[9][3] ),
    .ZN(_02932_));
 AOI22_X1 _07171_ (.A1(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[31][3] ),
    .A2(net96),
    .B1(net241),
    .B2(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[2][3] ),
    .ZN(_02933_));
 AOI22_X1 _07172_ (.A1(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[29][3] ),
    .A2(net143),
    .B1(net265),
    .B2(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[18][3] ),
    .ZN(_02934_));
 AOI21_X1 _07173_ (.A(net113),
    .B1(net75),
    .B2(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[28][3] ),
    .ZN(_02935_));
 NAND4_X1 _07174_ (.A1(_02932_),
    .A2(_02933_),
    .A3(_02934_),
    .A4(_02935_),
    .ZN(_02936_));
 AOI22_X1 _07175_ (.A1(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[5][3] ),
    .A2(net137),
    .B1(net205),
    .B2(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[13][3] ),
    .ZN(_02937_));
 AOI22_X1 _07176_ (.A1(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[15][3] ),
    .A2(net106),
    .B1(net271),
    .B2(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[12][3] ),
    .ZN(_02938_));
 AOI22_X1 _07177_ (.A1(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[16][3] ),
    .A2(net118),
    .B1(net91),
    .B2(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[10][3] ),
    .ZN(_02939_));
 AOI22_X1 _07178_ (.A1(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[17][3] ),
    .A2(net80),
    .B1(net82),
    .B2(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[21][3] ),
    .ZN(_02940_));
 NAND4_X1 _07179_ (.A1(_02937_),
    .A2(_02938_),
    .A3(_02939_),
    .A4(_02940_),
    .ZN(_02941_));
 AOI22_X1 _07180_ (.A1(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[23][3] ),
    .A2(net103),
    .B1(net169),
    .B2(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[26][3] ),
    .ZN(_02942_));
 AOI22_X1 _07181_ (.A1(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[20][3] ),
    .A2(net247),
    .B1(net235),
    .B2(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[11][3] ),
    .ZN(_02943_));
 AOI22_X1 _07182_ (.A1(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[8][3] ),
    .A2(net184),
    .B1(net125),
    .B2(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[4][3] ),
    .ZN(_02944_));
 AOI22_X2 _07183_ (.A1(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[7][3] ),
    .A2(net67),
    .B1(net210),
    .B2(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[30][3] ),
    .ZN(_02945_));
 NAND4_X2 _07184_ (.A1(_02942_),
    .A2(_02943_),
    .A3(_02944_),
    .A4(_02945_),
    .ZN(_02946_));
 NOR4_X2 _07185_ (.A1(_02931_),
    .A2(_02936_),
    .A3(_02941_),
    .A4(_02946_),
    .ZN(_02947_));
 OAI21_X1 _07186_ (.A(_01350_),
    .B1(net130),
    .B2(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[0][3] ),
    .ZN(_02948_));
 AOI22_X1 _07187_ (.A1(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[25][3] ),
    .A2(net154),
    .B1(net219),
    .B2(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[9][3] ),
    .ZN(_02949_));
 AOI22_X1 _07188_ (.A1(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[27][3] ),
    .A2(net189),
    .B1(net124),
    .B2(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[4][3] ),
    .ZN(_02950_));
 AOI22_X1 _07189_ (.A1(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[24][3] ),
    .A2(net74),
    .B1(net96),
    .B2(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[31][3] ),
    .ZN(_02951_));
 AOI22_X2 _07190_ (.A1(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[5][3] ),
    .A2(net137),
    .B1(net271),
    .B2(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[12][3] ),
    .ZN(_02952_));
 NAND4_X2 _07191_ (.A1(_02949_),
    .A2(_02950_),
    .A3(_02951_),
    .A4(_02952_),
    .ZN(_02953_));
 AOI22_X1 _07192_ (.A1(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[11][3] ),
    .A2(net234),
    .B1(net209),
    .B2(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[30][3] ),
    .ZN(_02954_));
 AOI22_X1 _07193_ (.A1(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[3][3] ),
    .A2(net64),
    .B1(net118),
    .B2(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[16][3] ),
    .ZN(_02955_));
 AOI22_X1 _07194_ (.A1(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[17][3] ),
    .A2(net80),
    .B1(net184),
    .B2(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[8][3] ),
    .ZN(_02956_));
 AOI21_X1 _07195_ (.A(net113),
    .B1(net259),
    .B2(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[1][3] ),
    .ZN(_02957_));
 NAND4_X1 _07196_ (.A1(_02954_),
    .A2(_02955_),
    .A3(_02956_),
    .A4(_02957_),
    .ZN(_02958_));
 AOI22_X1 _07197_ (.A1(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[28][3] ),
    .A2(net75),
    .B1(net241),
    .B2(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[2][3] ),
    .ZN(_02959_));
 AOI22_X1 _07198_ (.A1(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[23][3] ),
    .A2(net103),
    .B1(net169),
    .B2(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[26][3] ),
    .ZN(_02960_));
 AOI22_X1 _07199_ (.A1(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[6][3] ),
    .A2(net161),
    .B1(net67),
    .B2(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[7][3] ),
    .ZN(_02961_));
 AOI22_X1 _07200_ (.A1(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[29][3] ),
    .A2(net145),
    .B1(net247),
    .B2(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[20][3] ),
    .ZN(_02962_));
 NAND4_X1 _07201_ (.A1(_02959_),
    .A2(_02960_),
    .A3(_02961_),
    .A4(_02962_),
    .ZN(_02963_));
 AOI22_X1 _07202_ (.A1(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[10][3] ),
    .A2(net90),
    .B1(net85),
    .B2(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[14][3] ),
    .ZN(_02964_));
 AOI22_X1 _07203_ (.A1(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[13][3] ),
    .A2(net205),
    .B1(net195),
    .B2(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[19][3] ),
    .ZN(_02965_));
 AOI22_X1 _07204_ (.A1(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[15][3] ),
    .A2(net106),
    .B1(net224),
    .B2(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[22][3] ),
    .ZN(_02966_));
 AOI22_X1 _07205_ (.A1(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[18][3] ),
    .A2(net265),
    .B1(net82),
    .B2(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[21][3] ),
    .ZN(_02967_));
 NAND4_X1 _07206_ (.A1(_02964_),
    .A2(_02965_),
    .A3(_02966_),
    .A4(_02967_),
    .ZN(_02968_));
 NOR4_X2 _07207_ (.A1(_02953_),
    .A2(_02958_),
    .A3(_02963_),
    .A4(_02968_),
    .ZN(_02969_));
 OAI21_X1 _07208_ (.A(_01169_),
    .B1(net130),
    .B2(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[0][3] ),
    .ZN(_02970_));
 OAI22_X2 _07209_ (.A1(_02947_),
    .A2(_02948_),
    .B1(_02969_),
    .B2(_02970_),
    .ZN(_02971_));
 NOR4_X2 _07210_ (.A1(_02831_),
    .A2(_02879_),
    .A3(_02926_),
    .A4(_02971_),
    .ZN(_02972_));
 AOI22_X1 _07211_ (.A1(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[3][3] ),
    .A2(net64),
    .B1(net194),
    .B2(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[19][3] ),
    .ZN(_02973_));
 AOI22_X1 _07212_ (.A1(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[16][3] ),
    .A2(net116),
    .B1(net267),
    .B2(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[12][3] ),
    .ZN(_02974_));
 AOI22_X1 _07213_ (.A1(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[8][3] ),
    .A2(net179),
    .B1(net250),
    .B2(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[20][3] ),
    .ZN(_02975_));
 AOI22_X1 _07214_ (.A1(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[26][3] ),
    .A2(net173),
    .B1(net90),
    .B2(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[10][3] ),
    .ZN(_02976_));
 NAND4_X1 _07215_ (.A1(_02973_),
    .A2(_02974_),
    .A3(_02975_),
    .A4(_02976_),
    .ZN(_02977_));
 AOI22_X1 _07216_ (.A1(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[17][3] ),
    .A2(net79),
    .B1(net217),
    .B2(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[9][3] ),
    .ZN(_02978_));
 AOI22_X1 _07217_ (.A1(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[30][3] ),
    .A2(net208),
    .B1(net204),
    .B2(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[13][3] ),
    .ZN(_02979_));
 AOI22_X1 _07218_ (.A1(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[18][3] ),
    .A2(net263),
    .B1(net85),
    .B2(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[14][3] ),
    .ZN(_02980_));
 AOI21_X1 _07219_ (.A(net113),
    .B1(net100),
    .B2(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[23][3] ),
    .ZN(_02981_));
 NAND4_X1 _07220_ (.A1(_02978_),
    .A2(_02979_),
    .A3(_02980_),
    .A4(_02981_),
    .ZN(_02982_));
 AOI22_X1 _07221_ (.A1(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[15][3] ),
    .A2(net107),
    .B1(net131),
    .B2(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[5][3] ),
    .ZN(_02983_));
 AOI22_X1 _07222_ (.A1(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[25][3] ),
    .A2(net152),
    .B1(net255),
    .B2(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[1][3] ),
    .ZN(_02984_));
 AOI22_X1 _07223_ (.A1(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[29][3] ),
    .A2(net142),
    .B1(net233),
    .B2(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[11][3] ),
    .ZN(_02985_));
 AOI22_X1 _07224_ (.A1(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[7][3] ),
    .A2(net68),
    .B1(net93),
    .B2(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[31][3] ),
    .ZN(_02986_));
 NAND4_X1 _07225_ (.A1(_02983_),
    .A2(_02984_),
    .A3(_02985_),
    .A4(_02986_),
    .ZN(_02987_));
 AOI22_X1 _07226_ (.A1(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[4][3] ),
    .A2(net123),
    .B1(net82),
    .B2(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[21][3] ),
    .ZN(_02988_));
 AOI22_X1 _07227_ (.A1(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[27][3] ),
    .A2(net190),
    .B1(net226),
    .B2(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[22][3] ),
    .ZN(_02989_));
 AOI22_X1 _07228_ (.A1(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[28][3] ),
    .A2(net77),
    .B1(net162),
    .B2(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[6][3] ),
    .ZN(_02990_));
 AOI22_X1 _07229_ (.A1(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[24][3] ),
    .A2(net71),
    .B1(net240),
    .B2(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[2][3] ),
    .ZN(_02991_));
 NAND4_X1 _07230_ (.A1(_02988_),
    .A2(_02989_),
    .A3(_02990_),
    .A4(_02991_),
    .ZN(_02992_));
 OR4_X2 _07231_ (.A1(_02977_),
    .A2(_02982_),
    .A3(_02987_),
    .A4(_02992_),
    .ZN(_02993_));
 OAI21_X1 _07232_ (.A(_02993_),
    .B1(net130),
    .B2(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[0][3] ),
    .ZN(_02994_));
 AOI221_X2 _07233_ (.A(_00907_),
    .B1(_02781_),
    .B2(_02972_),
    .C1(_02994_),
    .C2(_01820_),
    .ZN(\rdata_o_n[3] ));
 OAI21_X1 _07234_ (.A(_01502_),
    .B1(_01064_),
    .B2(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[0][4] ),
    .ZN(_02995_));
 INV_X1 _07235_ (.A(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[19][4] ),
    .ZN(_02996_));
 INV_X1 _07236_ (.A(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[24][4] ),
    .ZN(_02997_));
 OAI33_X1 _07237_ (.A1(_02996_),
    .A2(_01015_),
    .A3(_00960_),
    .B1(_00954_),
    .B2(_00979_),
    .B3(_02997_),
    .ZN(_02998_));
 AOI221_X1 _07238_ (.A(_02998_),
    .B1(net89),
    .B2(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[10][4] ),
    .C1(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[17][4] ),
    .C2(net81),
    .ZN(_02999_));
 INV_X1 _07239_ (.A(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[8][4] ),
    .ZN(_03000_));
 NAND4_X4 _07240_ (.A1(_00953_),
    .A2(net10),
    .A3(_00946_),
    .A4(_00939_),
    .ZN(_03001_));
 INV_X1 _07241_ (.A(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[5][4] ),
    .ZN(_03002_));
 OAI22_X1 _07242_ (.A1(_03000_),
    .A2(_03001_),
    .B1(_02238_),
    .B2(_03002_),
    .ZN(_03003_));
 AOI221_X1 _07243_ (.A(_03003_),
    .B1(_01007_),
    .B2(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[13][4] ),
    .C1(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[14][4] ),
    .C2(net88),
    .ZN(_03004_));
 INV_X1 _07244_ (.A(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[27][4] ),
    .ZN(_03005_));
 INV_X1 _07245_ (.A(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[18][4] ),
    .ZN(_03006_));
 OAI22_X1 _07246_ (.A1(_03005_),
    .A2(_02555_),
    .B1(_02024_),
    .B2(_03006_),
    .ZN(_03007_));
 AOI221_X1 _07247_ (.A(_03007_),
    .B1(net70),
    .B2(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[7][4] ),
    .C1(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[22][4] ),
    .C2(_00996_),
    .ZN(_03008_));
 NAND2_X1 _07248_ (.A1(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[25][4] ),
    .A2(net151),
    .ZN(_03009_));
 NOR3_X4 _07249_ (.A1(_00953_),
    .A2(net10),
    .A3(_00946_),
    .ZN(_03010_));
 NAND3_X1 _07250_ (.A1(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[21][4] ),
    .A2(_01121_),
    .A3(_03010_),
    .ZN(_03011_));
 NAND2_X1 _07251_ (.A1(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[30][4] ),
    .A2(net215),
    .ZN(_03012_));
 NOR3_X4 _07252_ (.A1(net7),
    .A2(_00944_),
    .A3(_00946_),
    .ZN(_03013_));
 NAND3_X1 _07253_ (.A1(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[28][4] ),
    .A2(_01121_),
    .A3(_03013_),
    .ZN(_03014_));
 AND4_X1 _07254_ (.A1(_03009_),
    .A2(_03011_),
    .A3(_03012_),
    .A4(_03014_),
    .ZN(_03015_));
 AND4_X1 _07255_ (.A1(_02999_),
    .A2(_03004_),
    .A3(_03008_),
    .A4(_03015_),
    .ZN(_03016_));
 AOI22_X1 _07256_ (.A1(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[6][4] ),
    .A2(net156),
    .B1(net129),
    .B2(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[4][4] ),
    .ZN(_03017_));
 AOI22_X1 _07257_ (.A1(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[16][4] ),
    .A2(net121),
    .B1(net244),
    .B2(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[20][4] ),
    .ZN(_03018_));
 AOI22_X1 _07258_ (.A1(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[26][4] ),
    .A2(net167),
    .B1(net231),
    .B2(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[11][4] ),
    .ZN(_03019_));
 AOI22_X1 _07259_ (.A1(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[1][4] ),
    .A2(_00975_),
    .B1(_00989_),
    .B2(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[2][4] ),
    .ZN(_03020_));
 AND4_X1 _07260_ (.A1(_03017_),
    .A2(_03018_),
    .A3(_03019_),
    .A4(_03020_),
    .ZN(_03021_));
 AOI22_X1 _07261_ (.A1(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[31][4] ),
    .A2(_01149_),
    .B1(net274),
    .B2(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[12][4] ),
    .ZN(_03022_));
 AOI22_X1 _07262_ (.A1(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[3][4] ),
    .A2(net63),
    .B1(net112),
    .B2(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[15][4] ),
    .ZN(_03023_));
 INV_X1 _07263_ (.A(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[9][4] ),
    .ZN(_03024_));
 OAI21_X1 _07264_ (.A(_01064_),
    .B1(_01420_),
    .B2(_03024_),
    .ZN(_03025_));
 AOI221_X1 _07265_ (.A(_03025_),
    .B1(_01144_),
    .B2(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[23][4] ),
    .C1(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[29][4] ),
    .C2(_01050_),
    .ZN(_03026_));
 AND4_X1 _07266_ (.A1(_03021_),
    .A2(_03022_),
    .A3(_03023_),
    .A4(_03026_),
    .ZN(_03027_));
 AOI21_X1 _07267_ (.A(_02995_),
    .B1(_03016_),
    .B2(_03027_),
    .ZN(_03028_));
 OAI21_X1 _07268_ (.A(_00923_),
    .B1(_01064_),
    .B2(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[0][4] ),
    .ZN(_03029_));
 AOI22_X1 _07269_ (.A1(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[5][4] ),
    .A2(net136),
    .B1(net248),
    .B2(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[20][4] ),
    .ZN(_03030_));
 AOI22_X1 _07270_ (.A1(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[30][4] ),
    .A2(net207),
    .B1(net198),
    .B2(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[19][4] ),
    .ZN(_03031_));
 AOI22_X1 _07271_ (.A1(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[6][4] ),
    .A2(net160),
    .B1(net223),
    .B2(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[22][4] ),
    .ZN(_03032_));
 AOI22_X1 _07272_ (.A1(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[23][4] ),
    .A2(net98),
    .B1(net243),
    .B2(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[2][4] ),
    .ZN(_03033_));
 AND4_X1 _07273_ (.A1(_03030_),
    .A2(_03031_),
    .A3(_03032_),
    .A4(_03033_),
    .ZN(_03034_));
 AOI22_X1 _07274_ (.A1(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[17][4] ),
    .A2(net78),
    .B1(net65),
    .B2(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[3][4] ),
    .ZN(_03035_));
 AOI22_X1 _07275_ (.A1(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[7][4] ),
    .A2(net67),
    .B1(net91),
    .B2(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[10][4] ),
    .ZN(_03036_));
 INV_X1 _07276_ (.A(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[26][4] ),
    .ZN(_03037_));
 INV_X1 _07277_ (.A(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[12][4] ),
    .ZN(_03038_));
 OAI22_X1 _07278_ (.A1(_03037_),
    .A2(_01203_),
    .B1(_01426_),
    .B2(_03038_),
    .ZN(_03039_));
 AOI221_X1 _07279_ (.A(_03039_),
    .B1(net232),
    .B2(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[11][4] ),
    .C1(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[24][4] ),
    .C2(net72),
    .ZN(_03040_));
 AND4_X1 _07280_ (.A1(_03034_),
    .A2(_03035_),
    .A3(_03036_),
    .A4(_03040_),
    .ZN(_03041_));
 AOI22_X1 _07281_ (.A1(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[25][4] ),
    .A2(net149),
    .B1(_01149_),
    .B2(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[31][4] ),
    .ZN(_03042_));
 AOI22_X1 _07282_ (.A1(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[8][4] ),
    .A2(net182),
    .B1(net140),
    .B2(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[29][4] ),
    .ZN(_03043_));
 AND2_X1 _07283_ (.A1(_03042_),
    .A2(_03043_),
    .ZN(_03044_));
 AOI22_X1 _07284_ (.A1(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[27][4] ),
    .A2(net191),
    .B1(net206),
    .B2(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[13][4] ),
    .ZN(_03045_));
 AOI22_X1 _07285_ (.A1(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[16][4] ),
    .A2(net119),
    .B1(net128),
    .B2(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[4][4] ),
    .ZN(_03046_));
 AND2_X1 _07286_ (.A1(_03045_),
    .A2(_03046_),
    .ZN(_03047_));
 INV_X1 _07287_ (.A(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[21][4] ),
    .ZN(_03048_));
 INV_X1 _07288_ (.A(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[15][4] ),
    .ZN(_03049_));
 OAI33_X1 _07289_ (.A1(_03048_),
    .A2(_00979_),
    .A3(_00980_),
    .B1(_01005_),
    .B2(_00952_),
    .B3(_03049_),
    .ZN(_03050_));
 AOI221_X1 _07290_ (.A(_03050_),
    .B1(net258),
    .B2(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[1][4] ),
    .C1(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[18][4] ),
    .C2(net264),
    .ZN(_03051_));
 INV_X1 _07291_ (.A(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[9][4] ),
    .ZN(_03052_));
 OAI21_X1 _07292_ (.A(_01064_),
    .B1(_01420_),
    .B2(_03052_),
    .ZN(_03053_));
 AOI221_X1 _07293_ (.A(_03053_),
    .B1(net86),
    .B2(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[14][4] ),
    .C1(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[28][4] ),
    .C2(net75),
    .ZN(_03054_));
 AND4_X1 _07294_ (.A1(_03044_),
    .A2(_03047_),
    .A3(_03051_),
    .A4(_03054_),
    .ZN(_03055_));
 AOI21_X1 _07295_ (.A(_03029_),
    .B1(_03041_),
    .B2(_03055_),
    .ZN(_03056_));
 OR2_X1 _07296_ (.A1(_03028_),
    .A2(_03056_),
    .ZN(_03057_));
 AOI22_X1 _07297_ (.A1(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[23][4] ),
    .A2(net103),
    .B1(net265),
    .B2(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[18][4] ),
    .ZN(_03058_));
 AOI22_X1 _07298_ (.A1(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[15][4] ),
    .A2(net106),
    .B1(net169),
    .B2(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[26][4] ),
    .ZN(_03059_));
 AOI22_X1 _07299_ (.A1(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[8][4] ),
    .A2(net184),
    .B1(net205),
    .B2(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[13][4] ),
    .ZN(_03060_));
 AOI22_X2 _07300_ (.A1(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[3][4] ),
    .A2(net64),
    .B1(net235),
    .B2(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[11][4] ),
    .ZN(_03061_));
 NAND4_X2 _07301_ (.A1(_03058_),
    .A2(_03059_),
    .A3(_03060_),
    .A4(_03061_),
    .ZN(_03062_));
 AOI22_X1 _07302_ (.A1(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[12][4] ),
    .A2(net270),
    .B1(net220),
    .B2(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[9][4] ),
    .ZN(_03063_));
 AOI22_X1 _07303_ (.A1(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[24][4] ),
    .A2(net72),
    .B1(net85),
    .B2(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[14][4] ),
    .ZN(_03064_));
 AOI22_X1 _07304_ (.A1(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[28][4] ),
    .A2(net75),
    .B1(net259),
    .B2(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[1][4] ),
    .ZN(_03065_));
 AOI21_X1 _07305_ (.A(net113),
    .B1(net189),
    .B2(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[27][4] ),
    .ZN(_03066_));
 NAND4_X1 _07306_ (.A1(_03063_),
    .A2(_03064_),
    .A3(_03065_),
    .A4(_03066_),
    .ZN(_03067_));
 AOI22_X1 _07307_ (.A1(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[21][4] ),
    .A2(net82),
    .B1(net241),
    .B2(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[2][4] ),
    .ZN(_03068_));
 AOI22_X1 _07308_ (.A1(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[25][4] ),
    .A2(net155),
    .B1(net91),
    .B2(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[10][4] ),
    .ZN(_03069_));
 AOI22_X1 _07309_ (.A1(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[16][4] ),
    .A2(net118),
    .B1(net138),
    .B2(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[5][4] ),
    .ZN(_03070_));
 AOI22_X1 _07310_ (.A1(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[17][4] ),
    .A2(net80),
    .B1(net143),
    .B2(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[29][4] ),
    .ZN(_03071_));
 NAND4_X1 _07311_ (.A1(_03068_),
    .A2(_03069_),
    .A3(_03070_),
    .A4(_03071_),
    .ZN(_03072_));
 AOI22_X1 _07312_ (.A1(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[6][4] ),
    .A2(net164),
    .B1(_01009_),
    .B2(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[19][4] ),
    .ZN(_03073_));
 AOI22_X1 _07313_ (.A1(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[31][4] ),
    .A2(net96),
    .B1(net125),
    .B2(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[4][4] ),
    .ZN(_03074_));
 AOI22_X1 _07314_ (.A1(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[20][4] ),
    .A2(net247),
    .B1(net210),
    .B2(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[30][4] ),
    .ZN(_03075_));
 AOI22_X1 _07315_ (.A1(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[7][4] ),
    .A2(net67),
    .B1(net225),
    .B2(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[22][4] ),
    .ZN(_03076_));
 NAND4_X1 _07316_ (.A1(_03073_),
    .A2(_03074_),
    .A3(_03075_),
    .A4(_03076_),
    .ZN(_03077_));
 NOR4_X2 _07317_ (.A1(_03062_),
    .A2(_03067_),
    .A3(_03072_),
    .A4(_03077_),
    .ZN(_03078_));
 OAI21_X1 _07318_ (.A(_01350_),
    .B1(net130),
    .B2(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[0][4] ),
    .ZN(_03079_));
 OAI21_X1 _07319_ (.A(_01406_),
    .B1(_03078_),
    .B2(_03079_),
    .ZN(_03080_));
 INV_X1 _07320_ (.A(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[4][4] ),
    .ZN(_03081_));
 OAI21_X1 _07321_ (.A(_01064_),
    .B1(_00941_),
    .B2(_03081_),
    .ZN(_03082_));
 AOI221_X1 _07322_ (.A(_03082_),
    .B1(_00975_),
    .B2(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[1][4] ),
    .C1(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[24][4] ),
    .C2(net73),
    .ZN(_03083_));
 INV_X1 _07323_ (.A(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[29][4] ),
    .ZN(_03084_));
 INV_X1 _07324_ (.A(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[30][4] ),
    .ZN(_03085_));
 OAI22_X1 _07325_ (.A1(_03084_),
    .A2(_01425_),
    .B1(_01204_),
    .B2(_03085_),
    .ZN(_03086_));
 AOI221_X2 _07326_ (.A(_03086_),
    .B1(net156),
    .B2(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[6][4] ),
    .C1(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[10][4] ),
    .C2(net89),
    .ZN(_03087_));
 INV_X1 _07327_ (.A(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[21][4] ),
    .ZN(_03088_));
 INV_X1 _07328_ (.A(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[12][4] ),
    .ZN(_03089_));
 OAI33_X1 _07329_ (.A1(_03088_),
    .A2(_00979_),
    .A3(_00980_),
    .B1(_00970_),
    .B2(_00948_),
    .B3(_03089_),
    .ZN(_03090_));
 AOI221_X2 _07330_ (.A(_03090_),
    .B1(_01046_),
    .B2(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[25][4] ),
    .C1(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[27][4] ),
    .C2(_01021_),
    .ZN(_03091_));
 AOI22_X1 _07331_ (.A1(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[15][4] ),
    .A2(net112),
    .B1(net231),
    .B2(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[11][4] ),
    .ZN(_03092_));
 AOI22_X1 _07332_ (.A1(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[20][4] ),
    .A2(net244),
    .B1(net200),
    .B2(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[19][4] ),
    .ZN(_03093_));
 AND2_X1 _07333_ (.A1(_03092_),
    .A2(_03093_),
    .ZN(_03094_));
 NAND4_X2 _07334_ (.A1(_03083_),
    .A2(_03087_),
    .A3(_03091_),
    .A4(_03094_),
    .ZN(_03095_));
 AOI22_X1 _07335_ (.A1(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[5][4] ),
    .A2(net135),
    .B1(_00999_),
    .B2(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[9][4] ),
    .ZN(_03096_));
 AOI22_X1 _07336_ (.A1(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[3][4] ),
    .A2(net63),
    .B1(net206),
    .B2(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[13][4] ),
    .ZN(_03097_));
 AOI22_X1 _07337_ (.A1(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[16][4] ),
    .A2(net121),
    .B1(net264),
    .B2(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[18][4] ),
    .ZN(_03098_));
 AOI22_X2 _07338_ (.A1(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[7][4] ),
    .A2(net70),
    .B1(_00971_),
    .B2(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[14][4] ),
    .ZN(_03099_));
 NAND4_X2 _07339_ (.A1(_03096_),
    .A2(_03097_),
    .A3(_03098_),
    .A4(_03099_),
    .ZN(_03100_));
 AOI22_X1 _07340_ (.A1(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[26][4] ),
    .A2(net172),
    .B1(_01149_),
    .B2(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[31][4] ),
    .ZN(_03101_));
 AOI22_X1 _07341_ (.A1(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[23][4] ),
    .A2(_01144_),
    .B1(_00989_),
    .B2(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[2][4] ),
    .ZN(_03102_));
 AOI22_X1 _07342_ (.A1(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[28][4] ),
    .A2(_01032_),
    .B1(net176),
    .B2(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[8][4] ),
    .ZN(_03103_));
 AOI22_X2 _07343_ (.A1(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[17][4] ),
    .A2(net81),
    .B1(net228),
    .B2(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[22][4] ),
    .ZN(_03104_));
 NAND4_X2 _07344_ (.A1(_03101_),
    .A2(_03102_),
    .A3(_03103_),
    .A4(_03104_),
    .ZN(_03105_));
 NOR3_X4 _07345_ (.A1(_03095_),
    .A2(_03100_),
    .A3(_03105_),
    .ZN(_03106_));
 OAI21_X1 _07346_ (.A(_01731_),
    .B1(net130),
    .B2(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[0][4] ),
    .ZN(_03107_));
 AOI22_X1 _07347_ (.A1(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[16][4] ),
    .A2(net117),
    .B1(net153),
    .B2(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[25][4] ),
    .ZN(_03108_));
 AOI22_X1 _07348_ (.A1(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[31][4] ),
    .A2(net95),
    .B1(net194),
    .B2(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[19][4] ),
    .ZN(_03109_));
 AOI22_X1 _07349_ (.A1(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[23][4] ),
    .A2(net101),
    .B1(net251),
    .B2(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[20][4] ),
    .ZN(_03110_));
 AOI22_X1 _07350_ (.A1(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[26][4] ),
    .A2(net170),
    .B1(net234),
    .B2(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[11][4] ),
    .ZN(_03111_));
 NAND4_X1 _07351_ (.A1(_03108_),
    .A2(_03109_),
    .A3(_03110_),
    .A4(_03111_),
    .ZN(_03112_));
 AOI22_X1 _07352_ (.A1(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[8][4] ),
    .A2(net181),
    .B1(net68),
    .B2(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[7][4] ),
    .ZN(_03113_));
 AOI22_X1 _07353_ (.A1(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[15][4] ),
    .A2(net107),
    .B1(net204),
    .B2(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[13][4] ),
    .ZN(_03114_));
 MUX2_X1 _07354_ (.A(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[12][4] ),
    .B(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[14][4] ),
    .S(net8),
    .Z(_03115_));
 AOI221_X1 _07355_ (.A(net114),
    .B1(net92),
    .B2(_03115_),
    .C1(net242),
    .C2(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[2][4] ),
    .ZN(_03116_));
 NAND3_X1 _07356_ (.A1(_03113_),
    .A2(_03114_),
    .A3(_03116_),
    .ZN(_03117_));
 AOI22_X1 _07357_ (.A1(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[28][4] ),
    .A2(net77),
    .B1(net256),
    .B2(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[1][4] ),
    .ZN(_03118_));
 AOI22_X1 _07358_ (.A1(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[5][4] ),
    .A2(net132),
    .B1(net74),
    .B2(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[24][4] ),
    .ZN(_03119_));
 AOI22_X1 _07359_ (.A1(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[17][4] ),
    .A2(net80),
    .B1(net82),
    .B2(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[21][4] ),
    .ZN(_03120_));
 AOI22_X2 _07360_ (.A1(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[29][4] ),
    .A2(net142),
    .B1(net209),
    .B2(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[30][4] ),
    .ZN(_03121_));
 NAND4_X2 _07361_ (.A1(_03118_),
    .A2(_03119_),
    .A3(_03120_),
    .A4(_03121_),
    .ZN(_03122_));
 AOI22_X1 _07362_ (.A1(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[6][4] ),
    .A2(net163),
    .B1(net219),
    .B2(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[9][4] ),
    .ZN(_03123_));
 AOI22_X1 _07363_ (.A1(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[4][4] ),
    .A2(net124),
    .B1(net224),
    .B2(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[22][4] ),
    .ZN(_03124_));
 AOI22_X1 _07364_ (.A1(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[3][4] ),
    .A2(net64),
    .B1(net265),
    .B2(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[18][4] ),
    .ZN(_03125_));
 AOI22_X1 _07365_ (.A1(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[27][4] ),
    .A2(net190),
    .B1(net90),
    .B2(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[10][4] ),
    .ZN(_03126_));
 NAND4_X2 _07366_ (.A1(_03123_),
    .A2(_03124_),
    .A3(_03125_),
    .A4(_03126_),
    .ZN(_03127_));
 NOR4_X2 _07367_ (.A1(_03112_),
    .A2(_03117_),
    .A3(_03122_),
    .A4(_03127_),
    .ZN(_03128_));
 OAI21_X1 _07368_ (.A(_01539_),
    .B1(net130),
    .B2(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[0][4] ),
    .ZN(_03129_));
 OAI22_X1 _07369_ (.A1(_03106_),
    .A2(_03107_),
    .B1(_03128_),
    .B2(_03129_),
    .ZN(_03130_));
 AOI22_X1 _07370_ (.A1(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[11][4] ),
    .A2(net229),
    .B1(net213),
    .B2(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[30][4] ),
    .ZN(_03131_));
 AOI22_X1 _07371_ (.A1(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[12][4] ),
    .A2(_00950_),
    .B1(net238),
    .B2(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[2][4] ),
    .ZN(_03132_));
 AOI22_X1 _07372_ (.A1(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[17][4] ),
    .A2(net79),
    .B1(net218),
    .B2(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[9][4] ),
    .ZN(_03133_));
 AOI22_X1 _07373_ (.A1(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[15][4] ),
    .A2(net110),
    .B1(net88),
    .B2(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[14][4] ),
    .ZN(_03134_));
 NAND4_X2 _07374_ (.A1(_03131_),
    .A2(_03132_),
    .A3(_03133_),
    .A4(_03134_),
    .ZN(_03135_));
 AOI22_X1 _07375_ (.A1(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[28][4] ),
    .A2(net76),
    .B1(net131),
    .B2(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[5][4] ),
    .ZN(_03136_));
 AOI22_X1 _07376_ (.A1(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[23][4] ),
    .A2(net102),
    .B1(net126),
    .B2(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[4][4] ),
    .ZN(_03137_));
 AOI22_X1 _07377_ (.A1(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[8][4] ),
    .A2(net178),
    .B1(net254),
    .B2(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[1][4] ),
    .ZN(_03138_));
 AOI21_X1 _07378_ (.A(net114),
    .B1(net71),
    .B2(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[24][4] ),
    .ZN(_03139_));
 NAND4_X2 _07379_ (.A1(_03136_),
    .A2(_03137_),
    .A3(_03138_),
    .A4(_03139_),
    .ZN(_03140_));
 AOI22_X1 _07380_ (.A1(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[26][4] ),
    .A2(net174),
    .B1(net148),
    .B2(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[25][4] ),
    .ZN(_03141_));
 AOI22_X1 _07381_ (.A1(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[3][4] ),
    .A2(net66),
    .B1(net263),
    .B2(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[18][4] ),
    .ZN(_03142_));
 AOI22_X1 _07382_ (.A1(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[6][4] ),
    .A2(net158),
    .B1(net83),
    .B2(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[21][4] ),
    .ZN(_03143_));
 AOI22_X1 _07383_ (.A1(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[22][4] ),
    .A2(net222),
    .B1(net203),
    .B2(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[13][4] ),
    .ZN(_03144_));
 NAND4_X1 _07384_ (.A1(_03141_),
    .A2(_03142_),
    .A3(_03143_),
    .A4(_03144_),
    .ZN(_03145_));
 AOI22_X1 _07385_ (.A1(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[7][4] ),
    .A2(net69),
    .B1(net93),
    .B2(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[31][4] ),
    .ZN(_03146_));
 AOI22_X1 _07386_ (.A1(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[10][4] ),
    .A2(_00956_),
    .B1(net196),
    .B2(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[19][4] ),
    .ZN(_03147_));
 AOI22_X1 _07387_ (.A1(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[29][4] ),
    .A2(net144),
    .B1(net245),
    .B2(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[20][4] ),
    .ZN(_03148_));
 AOI22_X1 _07388_ (.A1(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[27][4] ),
    .A2(net188),
    .B1(net120),
    .B2(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[16][4] ),
    .ZN(_03149_));
 NAND4_X1 _07389_ (.A1(_03146_),
    .A2(_03147_),
    .A3(_03148_),
    .A4(_03149_),
    .ZN(_03150_));
 NOR4_X2 _07390_ (.A1(_03135_),
    .A2(_03140_),
    .A3(_03145_),
    .A4(_03150_),
    .ZN(_03151_));
 OAI21_X1 _07391_ (.A(_01295_),
    .B1(net130),
    .B2(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[0][4] ),
    .ZN(_03152_));
 AOI22_X1 _07392_ (.A1(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[1][4] ),
    .A2(net253),
    .B1(net206),
    .B2(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[13][4] ),
    .ZN(_03153_));
 AOI22_X1 _07393_ (.A1(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[20][4] ),
    .A2(net252),
    .B1(net237),
    .B2(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[11][4] ),
    .ZN(_03154_));
 AOI22_X1 _07394_ (.A1(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[14][4] ),
    .A2(net87),
    .B1(_00999_),
    .B2(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[9][4] ),
    .ZN(_03155_));
 AOI22_X1 _07395_ (.A1(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[12][4] ),
    .A2(net272),
    .B1(net211),
    .B2(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[30][4] ),
    .ZN(_03156_));
 NAND4_X1 _07396_ (.A1(_03153_),
    .A2(_03154_),
    .A3(_03155_),
    .A4(_03156_),
    .ZN(_03157_));
 AOI22_X1 _07397_ (.A1(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[31][4] ),
    .A2(_01149_),
    .B1(net243),
    .B2(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[2][4] ),
    .ZN(_03158_));
 AOI22_X1 _07398_ (.A1(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[3][4] ),
    .A2(net65),
    .B1(net139),
    .B2(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[5][4] ),
    .ZN(_03159_));
 AOI22_X1 _07399_ (.A1(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[15][4] ),
    .A2(net109),
    .B1(net225),
    .B2(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[22][4] ),
    .ZN(_03160_));
 AOI21_X1 _07400_ (.A(_01119_),
    .B1(net182),
    .B2(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[8][4] ),
    .ZN(_03161_));
 NAND4_X2 _07401_ (.A1(_03158_),
    .A2(_03159_),
    .A3(_03160_),
    .A4(_03161_),
    .ZN(_03162_));
 AOI22_X1 _07402_ (.A1(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[26][4] ),
    .A2(net171),
    .B1(net128),
    .B2(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[4][4] ),
    .ZN(_03163_));
 AOI22_X1 _07403_ (.A1(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[28][4] ),
    .A2(_01032_),
    .B1(net198),
    .B2(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[19][4] ),
    .ZN(_03164_));
 AOI22_X1 _07404_ (.A1(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[10][4] ),
    .A2(net89),
    .B1(net264),
    .B2(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[18][4] ),
    .ZN(_03165_));
 AOI22_X2 _07405_ (.A1(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[16][4] ),
    .A2(net119),
    .B1(net84),
    .B2(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[21][4] ),
    .ZN(_03166_));
 NAND4_X2 _07406_ (.A1(_03163_),
    .A2(_03164_),
    .A3(_03165_),
    .A4(_03166_),
    .ZN(_03167_));
 AOI22_X1 _07407_ (.A1(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[17][4] ),
    .A2(net78),
    .B1(net192),
    .B2(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[27][4] ),
    .ZN(_03168_));
 AOI22_X1 _07408_ (.A1(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[29][4] ),
    .A2(net140),
    .B1(net73),
    .B2(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[24][4] ),
    .ZN(_03169_));
 AOI22_X1 _07409_ (.A1(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[25][4] ),
    .A2(net149),
    .B1(_01076_),
    .B2(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[7][4] ),
    .ZN(_03170_));
 AOI22_X1 _07410_ (.A1(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[23][4] ),
    .A2(net99),
    .B1(net160),
    .B2(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[6][4] ),
    .ZN(_03171_));
 NAND4_X1 _07411_ (.A1(_03168_),
    .A2(_03169_),
    .A3(_03170_),
    .A4(_03171_),
    .ZN(_03172_));
 NOR4_X2 _07412_ (.A1(_03157_),
    .A2(_03162_),
    .A3(_03167_),
    .A4(_03172_),
    .ZN(_03173_));
 OAI21_X1 _07413_ (.A(_01408_),
    .B1(net130),
    .B2(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[0][4] ),
    .ZN(_03174_));
 OAI22_X2 _07414_ (.A1(_03151_),
    .A2(_03152_),
    .B1(_03173_),
    .B2(_03174_),
    .ZN(_03175_));
 NOR4_X1 _07415_ (.A1(_03057_),
    .A2(_03080_),
    .A3(_03130_),
    .A4(_03175_),
    .ZN(_03176_));
 AOI22_X1 _07416_ (.A1(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[17][4] ),
    .A2(net80),
    .B1(net126),
    .B2(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[4][4] ),
    .ZN(_03177_));
 AOI22_X1 _07417_ (.A1(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[28][4] ),
    .A2(net77),
    .B1(net68),
    .B2(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[7][4] ),
    .ZN(_03178_));
 AOI22_X1 _07418_ (.A1(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[25][4] ),
    .A2(net152),
    .B1(net87),
    .B2(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[14][4] ),
    .ZN(_03179_));
 AOI22_X1 _07419_ (.A1(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[6][4] ),
    .A2(net164),
    .B1(net212),
    .B2(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[30][4] ),
    .ZN(_03180_));
 NAND4_X1 _07420_ (.A1(_03177_),
    .A2(_03178_),
    .A3(_03179_),
    .A4(_03180_),
    .ZN(_03181_));
 AOI22_X1 _07421_ (.A1(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[15][4] ),
    .A2(net108),
    .B1(net218),
    .B2(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[9][4] ),
    .ZN(_03182_));
 AOI22_X1 _07422_ (.A1(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[27][4] ),
    .A2(net188),
    .B1(net242),
    .B2(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[2][4] ),
    .ZN(_03183_));
 AOI22_X1 _07423_ (.A1(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[12][4] ),
    .A2(net269),
    .B1(net83),
    .B2(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[21][4] ),
    .ZN(_03184_));
 AOI21_X1 _07424_ (.A(net114),
    .B1(net226),
    .B2(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[22][4] ),
    .ZN(_03185_));
 NAND4_X1 _07425_ (.A1(_03182_),
    .A2(_03183_),
    .A3(_03184_),
    .A4(_03185_),
    .ZN(_03186_));
 AOI22_X1 _07426_ (.A1(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[8][4] ),
    .A2(net180),
    .B1(net236),
    .B2(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[11][4] ),
    .ZN(_03187_));
 AOI22_X1 _07427_ (.A1(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[16][4] ),
    .A2(net116),
    .B1(net263),
    .B2(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[18][4] ),
    .ZN(_03188_));
 AOI22_X1 _07428_ (.A1(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[5][4] ),
    .A2(net132),
    .B1(net203),
    .B2(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[13][4] ),
    .ZN(_03189_));
 AOI22_X1 _07429_ (.A1(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[26][4] ),
    .A2(net173),
    .B1(net193),
    .B2(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[19][4] ),
    .ZN(_03190_));
 NAND4_X1 _07430_ (.A1(_03187_),
    .A2(_03188_),
    .A3(_03189_),
    .A4(_03190_),
    .ZN(_03191_));
 AOI22_X1 _07431_ (.A1(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[31][4] ),
    .A2(net95),
    .B1(net90),
    .B2(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[10][4] ),
    .ZN(_03192_));
 AOI22_X1 _07432_ (.A1(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[23][4] ),
    .A2(net101),
    .B1(net260),
    .B2(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[1][4] ),
    .ZN(_03193_));
 AOI22_X1 _07433_ (.A1(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[3][4] ),
    .A2(net64),
    .B1(net74),
    .B2(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[24][4] ),
    .ZN(_03194_));
 AOI22_X1 _07434_ (.A1(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[29][4] ),
    .A2(net144),
    .B1(net251),
    .B2(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[20][4] ),
    .ZN(_03195_));
 NAND4_X1 _07435_ (.A1(_03192_),
    .A2(_03193_),
    .A3(_03194_),
    .A4(_03195_),
    .ZN(_03196_));
 NOR4_X1 _07436_ (.A1(_03181_),
    .A2(_03186_),
    .A3(_03191_),
    .A4(_03196_),
    .ZN(_03197_));
 OAI21_X1 _07437_ (.A(_01700_),
    .B1(net130),
    .B2(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[0][4] ),
    .ZN(_03198_));
 AOI22_X1 _07438_ (.A1(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[5][4] ),
    .A2(net135),
    .B1(net200),
    .B2(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[19][4] ),
    .ZN(_03199_));
 AOI22_X1 _07439_ (.A1(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[29][4] ),
    .A2(net141),
    .B1(net262),
    .B2(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[1][4] ),
    .ZN(_03200_));
 AOI22_X1 _07440_ (.A1(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[24][4] ),
    .A2(_01059_),
    .B1(net246),
    .B2(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[20][4] ),
    .ZN(_03201_));
 AOI22_X1 _07441_ (.A1(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[15][4] ),
    .A2(net111),
    .B1(net227),
    .B2(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[22][4] ),
    .ZN(_03202_));
 NAND4_X1 _07442_ (.A1(_03199_),
    .A2(_03200_),
    .A3(_03201_),
    .A4(_03202_),
    .ZN(_03203_));
 AOI22_X2 _07443_ (.A1(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[14][4] ),
    .A2(net88),
    .B1(net221),
    .B2(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[9][4] ),
    .ZN(_03204_));
 AOI22_X1 _07444_ (.A1(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[17][4] ),
    .A2(net81),
    .B1(net167),
    .B2(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[26][4] ),
    .ZN(_03205_));
 AOI22_X1 _07445_ (.A1(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[28][4] ),
    .A2(_01032_),
    .B1(_00981_),
    .B2(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[21][4] ),
    .ZN(_03206_));
 AOI21_X1 _07446_ (.A(net115),
    .B1(net63),
    .B2(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[3][4] ),
    .ZN(_03207_));
 NAND4_X2 _07447_ (.A1(_03204_),
    .A2(_03205_),
    .A3(_03206_),
    .A4(_03207_),
    .ZN(_03208_));
 AOI22_X1 _07448_ (.A1(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[8][4] ),
    .A2(net177),
    .B1(net239),
    .B2(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[2][4] ),
    .ZN(_03209_));
 AOI22_X1 _07449_ (.A1(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[23][4] ),
    .A2(net97),
    .B1(net216),
    .B2(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[30][4] ),
    .ZN(_03210_));
 AOI22_X1 _07450_ (.A1(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[16][4] ),
    .A2(net122),
    .B1(_00964_),
    .B2(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[18][4] ),
    .ZN(_03211_));
 AOI22_X2 _07451_ (.A1(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[27][4] ),
    .A2(net186),
    .B1(net70),
    .B2(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[7][4] ),
    .ZN(_03212_));
 NAND4_X2 _07452_ (.A1(_03209_),
    .A2(_03210_),
    .A3(_03211_),
    .A4(_03212_),
    .ZN(_03213_));
 AOI22_X1 _07453_ (.A1(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[31][4] ),
    .A2(net94),
    .B1(_01007_),
    .B2(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[13][4] ),
    .ZN(_03214_));
 AOI22_X2 _07454_ (.A1(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[25][4] ),
    .A2(net151),
    .B1(net273),
    .B2(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[12][4] ),
    .ZN(_03215_));
 AOI22_X1 _07455_ (.A1(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[6][4] ),
    .A2(net159),
    .B1(net129),
    .B2(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[4][4] ),
    .ZN(_03216_));
 AOI22_X2 _07456_ (.A1(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[10][4] ),
    .A2(net89),
    .B1(_00993_),
    .B2(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[11][4] ),
    .ZN(_03217_));
 NAND4_X2 _07457_ (.A1(_03214_),
    .A2(_03215_),
    .A3(_03216_),
    .A4(_03217_),
    .ZN(_03218_));
 NOR4_X2 _07458_ (.A1(_03203_),
    .A2(_03208_),
    .A3(_03213_),
    .A4(_03218_),
    .ZN(_03219_));
 OAI21_X1 _07459_ (.A(_01662_),
    .B1(net130),
    .B2(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[0][4] ),
    .ZN(_03220_));
 OAI22_X1 _07460_ (.A1(_03197_),
    .A2(_03198_),
    .B1(_03219_),
    .B2(_03220_),
    .ZN(_03221_));
 AOI22_X1 _07461_ (.A1(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[21][4] ),
    .A2(net83),
    .B1(net238),
    .B2(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[2][4] ),
    .ZN(_03222_));
 AOI22_X1 _07462_ (.A1(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[28][4] ),
    .A2(net76),
    .B1(net246),
    .B2(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[20][4] ),
    .ZN(_03223_));
 AOI22_X1 _07463_ (.A1(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[6][4] ),
    .A2(net157),
    .B1(net126),
    .B2(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[4][4] ),
    .ZN(_03224_));
 AOI22_X1 _07464_ (.A1(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[7][4] ),
    .A2(net69),
    .B1(net229),
    .B2(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[11][4] ),
    .ZN(_03225_));
 NAND4_X2 _07465_ (.A1(_03222_),
    .A2(_03223_),
    .A3(_03224_),
    .A4(_03225_),
    .ZN(_03226_));
 AOI22_X1 _07466_ (.A1(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[3][4] ),
    .A2(_01102_),
    .B1(net147),
    .B2(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[25][4] ),
    .ZN(_03227_));
 AOI22_X1 _07467_ (.A1(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[5][4] ),
    .A2(net133),
    .B1(net218),
    .B2(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[9][4] ),
    .ZN(_03228_));
 MUX2_X1 _07468_ (.A(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[24][4] ),
    .B(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[26][4] ),
    .S(net8),
    .Z(_03229_));
 AOI22_X1 _07469_ (.A1(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[8][4] ),
    .A2(_00939_),
    .B1(_03229_),
    .B2(net1),
    .ZN(_03230_));
 INV_X1 _07470_ (.A(_03230_),
    .ZN(_03231_));
 AOI221_X2 _07471_ (.A(net115),
    .B1(net199),
    .B2(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[19][4] ),
    .C1(_03231_),
    .C2(_02912_),
    .ZN(_03232_));
 NAND3_X2 _07472_ (.A1(_03227_),
    .A2(_03228_),
    .A3(_03232_),
    .ZN(_03233_));
 AOI22_X1 _07473_ (.A1(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[15][4] ),
    .A2(net110),
    .B1(net94),
    .B2(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[31][4] ),
    .ZN(_03234_));
 AOI22_X1 _07474_ (.A1(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[12][4] ),
    .A2(net273),
    .B1(_00964_),
    .B2(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[18][4] ),
    .ZN(_03235_));
 AOI22_X1 _07475_ (.A1(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[27][4] ),
    .A2(net187),
    .B1(net203),
    .B2(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[13][4] ),
    .ZN(_03236_));
 AOI22_X1 _07476_ (.A1(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[10][4] ),
    .A2(net89),
    .B1(net88),
    .B2(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[14][4] ),
    .ZN(_03237_));
 NAND4_X2 _07477_ (.A1(_03234_),
    .A2(_03235_),
    .A3(_03236_),
    .A4(_03237_),
    .ZN(_03238_));
 AOI222_X2 _07478_ (.A1(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[23][4] ),
    .A2(net102),
    .B1(net120),
    .B2(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[16][4] ),
    .C1(net227),
    .C2(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[22][4] ),
    .ZN(_03239_));
 AOI22_X1 _07479_ (.A1(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[17][4] ),
    .A2(net79),
    .B1(net261),
    .B2(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[1][4] ),
    .ZN(_03240_));
 AOI22_X1 _07480_ (.A1(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[29][4] ),
    .A2(net141),
    .B1(net213),
    .B2(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[30][4] ),
    .ZN(_03241_));
 NAND3_X2 _07481_ (.A1(_03239_),
    .A2(_03240_),
    .A3(_03241_),
    .ZN(_03242_));
 NOR4_X4 _07482_ (.A1(_03226_),
    .A2(_03233_),
    .A3(_03238_),
    .A4(_03242_),
    .ZN(_03243_));
 OAI21_X1 _07483_ (.A(_01583_),
    .B1(net130),
    .B2(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[0][4] ),
    .ZN(_03244_));
 AOI22_X1 _07484_ (.A1(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[7][4] ),
    .A2(net68),
    .B1(net263),
    .B2(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[18][4] ),
    .ZN(_03245_));
 AOI22_X1 _07485_ (.A1(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[28][4] ),
    .A2(net76),
    .B1(net222),
    .B2(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[22][4] ),
    .ZN(_03246_));
 AOI22_X1 _07486_ (.A1(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[25][4] ),
    .A2(net152),
    .B1(net208),
    .B2(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[30][4] ),
    .ZN(_03247_));
 AOI22_X1 _07487_ (.A1(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[3][4] ),
    .A2(net66),
    .B1(net108),
    .B2(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[15][4] ),
    .ZN(_03248_));
 NAND4_X1 _07488_ (.A1(_03245_),
    .A2(_03246_),
    .A3(_03247_),
    .A4(_03248_),
    .ZN(_03249_));
 AOI22_X1 _07489_ (.A1(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[8][4] ),
    .A2(net180),
    .B1(net193),
    .B2(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[19][4] ),
    .ZN(_03250_));
 AOI22_X1 _07490_ (.A1(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[23][4] ),
    .A2(net100),
    .B1(net233),
    .B2(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[11][4] ),
    .ZN(_03251_));
 MUX2_X1 _07491_ (.A(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[12][4] ),
    .B(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[14][4] ),
    .S(net8),
    .Z(_03252_));
 AOI221_X1 _07492_ (.A(net114),
    .B1(net92),
    .B2(_03252_),
    .C1(net254),
    .C2(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[1][4] ),
    .ZN(_03253_));
 NAND3_X1 _07493_ (.A1(_03250_),
    .A2(_03251_),
    .A3(_03253_),
    .ZN(_03254_));
 AOI22_X1 _07494_ (.A1(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[5][4] ),
    .A2(net131),
    .B1(net240),
    .B2(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[2][4] ),
    .ZN(_03255_));
 AOI22_X1 _07495_ (.A1(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[29][4] ),
    .A2(net144),
    .B1(net71),
    .B2(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[24][4] ),
    .ZN(_03256_));
 AOI22_X1 _07496_ (.A1(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[20][4] ),
    .A2(net250),
    .B1(net217),
    .B2(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[9][4] ),
    .ZN(_03257_));
 AOI22_X2 _07497_ (.A1(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[27][4] ),
    .A2(net188),
    .B1(net116),
    .B2(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[16][4] ),
    .ZN(_03258_));
 NAND4_X2 _07498_ (.A1(_03255_),
    .A2(_03256_),
    .A3(_03257_),
    .A4(_03258_),
    .ZN(_03259_));
 AOI22_X1 _07499_ (.A1(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[17][4] ),
    .A2(net79),
    .B1(net123),
    .B2(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[4][4] ),
    .ZN(_03260_));
 AOI22_X1 _07500_ (.A1(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[31][4] ),
    .A2(net93),
    .B1(net83),
    .B2(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[21][4] ),
    .ZN(_03261_));
 AOI22_X1 _07501_ (.A1(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[6][4] ),
    .A2(net162),
    .B1(net204),
    .B2(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[13][4] ),
    .ZN(_03262_));
 AOI22_X1 _07502_ (.A1(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[26][4] ),
    .A2(net175),
    .B1(net90),
    .B2(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[10][4] ),
    .ZN(_03263_));
 NAND4_X1 _07503_ (.A1(_03260_),
    .A2(_03261_),
    .A3(_03262_),
    .A4(_03263_),
    .ZN(_03264_));
 NOR4_X2 _07504_ (.A1(_03249_),
    .A2(_03254_),
    .A3(_03259_),
    .A4(_03264_),
    .ZN(_03265_));
 OAI21_X1 _07505_ (.A(_01401_),
    .B1(net130),
    .B2(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[0][4] ),
    .ZN(_03266_));
 OAI22_X2 _07506_ (.A1(_03243_),
    .A2(_03244_),
    .B1(_03265_),
    .B2(_03266_),
    .ZN(_03267_));
 AOI22_X1 _07507_ (.A1(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[25][4] ),
    .A2(net154),
    .B1(net124),
    .B2(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[4][4] ),
    .ZN(_03268_));
 AOI22_X1 _07508_ (.A1(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[16][4] ),
    .A2(net118),
    .B1(net169),
    .B2(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[26][4] ),
    .ZN(_03269_));
 AOI22_X1 _07509_ (.A1(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[6][4] ),
    .A2(net161),
    .B1(net82),
    .B2(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[21][4] ),
    .ZN(_03270_));
 AOI22_X2 _07510_ (.A1(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[23][4] ),
    .A2(net103),
    .B1(net219),
    .B2(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[9][4] ),
    .ZN(_03271_));
 NAND4_X2 _07511_ (.A1(_03268_),
    .A2(_03269_),
    .A3(_03270_),
    .A4(_03271_),
    .ZN(_03272_));
 AOI22_X1 _07512_ (.A1(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[10][4] ),
    .A2(net90),
    .B1(net85),
    .B2(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[14][4] ),
    .ZN(_03273_));
 AOI22_X1 _07513_ (.A1(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[15][4] ),
    .A2(net106),
    .B1(net234),
    .B2(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[11][4] ),
    .ZN(_03274_));
 AOI22_X1 _07514_ (.A1(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[24][4] ),
    .A2(net74),
    .B1(net241),
    .B2(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[2][4] ),
    .ZN(_03275_));
 AOI21_X1 _07515_ (.A(net113),
    .B1(net209),
    .B2(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[30][4] ),
    .ZN(_03276_));
 NAND4_X1 _07516_ (.A1(_03273_),
    .A2(_03274_),
    .A3(_03275_),
    .A4(_03276_),
    .ZN(_03277_));
 AOI22_X1 _07517_ (.A1(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[17][4] ),
    .A2(net80),
    .B1(net145),
    .B2(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[29][4] ),
    .ZN(_03278_));
 AOI22_X1 _07518_ (.A1(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[27][4] ),
    .A2(net189),
    .B1(net75),
    .B2(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[28][4] ),
    .ZN(_03279_));
 AOI22_X1 _07519_ (.A1(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[5][4] ),
    .A2(net137),
    .B1(net67),
    .B2(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[7][4] ),
    .ZN(_03280_));
 AOI22_X2 _07520_ (.A1(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[1][4] ),
    .A2(net259),
    .B1(net205),
    .B2(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[13][4] ),
    .ZN(_03281_));
 NAND4_X2 _07521_ (.A1(_03278_),
    .A2(_03279_),
    .A3(_03280_),
    .A4(_03281_),
    .ZN(_03282_));
 AOI22_X1 _07522_ (.A1(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[8][4] ),
    .A2(net184),
    .B1(net96),
    .B2(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[31][4] ),
    .ZN(_03283_));
 AOI22_X1 _07523_ (.A1(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[18][4] ),
    .A2(net265),
    .B1(net249),
    .B2(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[20][4] ),
    .ZN(_03284_));
 AOI22_X1 _07524_ (.A1(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[12][4] ),
    .A2(net271),
    .B1(net195),
    .B2(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[19][4] ),
    .ZN(_03285_));
 AOI22_X1 _07525_ (.A1(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[3][4] ),
    .A2(net64),
    .B1(net224),
    .B2(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[22][4] ),
    .ZN(_03286_));
 NAND4_X1 _07526_ (.A1(_03283_),
    .A2(_03284_),
    .A3(_03285_),
    .A4(_03286_),
    .ZN(_03287_));
 NOR4_X2 _07527_ (.A1(_03272_),
    .A2(_03277_),
    .A3(_03282_),
    .A4(_03287_),
    .ZN(_03288_));
 OAI21_X1 _07528_ (.A(_01169_),
    .B1(net130),
    .B2(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[0][4] ),
    .ZN(_03289_));
 AOI22_X1 _07529_ (.A1(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[23][4] ),
    .A2(net97),
    .B1(net159),
    .B2(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[6][4] ),
    .ZN(_03290_));
 AOI22_X1 _07530_ (.A1(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[28][4] ),
    .A2(net76),
    .B1(net227),
    .B2(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[22][4] ),
    .ZN(_03291_));
 AOI22_X2 _07531_ (.A1(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[4][4] ),
    .A2(net127),
    .B1(net273),
    .B2(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[12][4] ),
    .ZN(_03292_));
 AOI22_X2 _07532_ (.A1(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[17][4] ),
    .A2(net81),
    .B1(net63),
    .B2(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[3][4] ),
    .ZN(_03293_));
 NAND4_X2 _07533_ (.A1(_03290_),
    .A2(_03291_),
    .A3(_03292_),
    .A4(_03293_),
    .ZN(_03294_));
 AOI22_X1 _07534_ (.A1(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[25][4] ),
    .A2(net147),
    .B1(net216),
    .B2(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[30][4] ),
    .ZN(_03295_));
 AOI22_X1 _07535_ (.A1(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[24][4] ),
    .A2(_01059_),
    .B1(_00981_),
    .B2(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[21][4] ),
    .ZN(_03296_));
 AOI22_X1 _07536_ (.A1(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[8][4] ),
    .A2(net185),
    .B1(net133),
    .B2(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[5][4] ),
    .ZN(_03297_));
 AOI21_X1 _07537_ (.A(net115),
    .B1(net202),
    .B2(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[19][4] ),
    .ZN(_03298_));
 NAND4_X2 _07538_ (.A1(_03295_),
    .A2(_03296_),
    .A3(_03297_),
    .A4(_03298_),
    .ZN(_03299_));
 AOI22_X1 _07539_ (.A1(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[27][4] ),
    .A2(net187),
    .B1(net166),
    .B2(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[26][4] ),
    .ZN(_03300_));
 AOI22_X2 _07540_ (.A1(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[7][4] ),
    .A2(net70),
    .B1(_00964_),
    .B2(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[18][4] ),
    .ZN(_03301_));
 AOI22_X1 _07541_ (.A1(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[29][4] ),
    .A2(net141),
    .B1(net218),
    .B2(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[9][4] ),
    .ZN(_03302_));
 AOI22_X2 _07542_ (.A1(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[15][4] ),
    .A2(net110),
    .B1(net94),
    .B2(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[31][4] ),
    .ZN(_03303_));
 NAND4_X2 _07543_ (.A1(_03300_),
    .A2(_03301_),
    .A3(_03302_),
    .A4(_03303_),
    .ZN(_03304_));
 AOI22_X1 _07544_ (.A1(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[16][4] ),
    .A2(net122),
    .B1(net261),
    .B2(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[1][4] ),
    .ZN(_03305_));
 AOI22_X1 _07545_ (.A1(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[14][4] ),
    .A2(net88),
    .B1(net239),
    .B2(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[2][4] ),
    .ZN(_03306_));
 AOI22_X1 _07546_ (.A1(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[10][4] ),
    .A2(net89),
    .B1(net230),
    .B2(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[11][4] ),
    .ZN(_03307_));
 AOI22_X2 _07547_ (.A1(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[20][4] ),
    .A2(net246),
    .B1(net203),
    .B2(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[13][4] ),
    .ZN(_03308_));
 NAND4_X2 _07548_ (.A1(_03305_),
    .A2(_03306_),
    .A3(_03307_),
    .A4(_03308_),
    .ZN(_03309_));
 NOR4_X4 _07549_ (.A1(_03294_),
    .A2(_03299_),
    .A3(_03304_),
    .A4(_03309_),
    .ZN(_03310_));
 OAI21_X1 _07550_ (.A(_01623_),
    .B1(net130),
    .B2(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[0][4] ),
    .ZN(_03311_));
 OAI22_X1 _07551_ (.A1(_03288_),
    .A2(_03289_),
    .B1(_03310_),
    .B2(_03311_),
    .ZN(_03312_));
 AOI22_X1 _07552_ (.A1(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[3][4] ),
    .A2(net65),
    .B1(_01097_),
    .B2(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[16][4] ),
    .ZN(_03313_));
 AOI22_X1 _07553_ (.A1(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[31][4] ),
    .A2(net96),
    .B1(net220),
    .B2(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[9][4] ),
    .ZN(_03314_));
 AOI22_X1 _07554_ (.A1(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[25][4] ),
    .A2(net155),
    .B1(net125),
    .B2(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[4][4] ),
    .ZN(_03315_));
 AOI22_X1 _07555_ (.A1(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[23][4] ),
    .A2(net105),
    .B1(net83),
    .B2(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[21][4] ),
    .ZN(_03316_));
 NAND4_X1 _07556_ (.A1(_03313_),
    .A2(_03314_),
    .A3(_03315_),
    .A4(_03316_),
    .ZN(_03317_));
 AOI22_X1 _07557_ (.A1(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[26][4] ),
    .A2(net168),
    .B1(net205),
    .B2(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[13][4] ),
    .ZN(_03318_));
 AOI22_X1 _07558_ (.A1(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[10][4] ),
    .A2(net91),
    .B1(net86),
    .B2(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[14][4] ),
    .ZN(_03319_));
 AOI22_X1 _07559_ (.A1(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[17][4] ),
    .A2(net78),
    .B1(net191),
    .B2(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[27][4] ),
    .ZN(_03320_));
 AOI21_X1 _07560_ (.A(net113),
    .B1(net138),
    .B2(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[5][4] ),
    .ZN(_03321_));
 NAND4_X1 _07561_ (.A1(_03318_),
    .A2(_03319_),
    .A3(_03320_),
    .A4(_03321_),
    .ZN(_03322_));
 AOI22_X1 _07562_ (.A1(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[20][4] ),
    .A2(net249),
    .B1(net212),
    .B2(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[30][4] ),
    .ZN(_03323_));
 AOI22_X1 _07563_ (.A1(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[29][4] ),
    .A2(net145),
    .B1(net235),
    .B2(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[11][4] ),
    .ZN(_03324_));
 AOI22_X1 _07564_ (.A1(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[8][4] ),
    .A2(_01034_),
    .B1(net265),
    .B2(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[18][4] ),
    .ZN(_03325_));
 AOI22_X1 _07565_ (.A1(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[15][4] ),
    .A2(net108),
    .B1(net271),
    .B2(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[12][4] ),
    .ZN(_03326_));
 NAND4_X1 _07566_ (.A1(_03323_),
    .A2(_03324_),
    .A3(_03325_),
    .A4(_03326_),
    .ZN(_03327_));
 AOI22_X1 _07567_ (.A1(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[7][4] ),
    .A2(net68),
    .B1(_01009_),
    .B2(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[19][4] ),
    .ZN(_03328_));
 AOI22_X1 _07568_ (.A1(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[28][4] ),
    .A2(net75),
    .B1(net258),
    .B2(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[1][4] ),
    .ZN(_03329_));
 AOI22_X1 _07569_ (.A1(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[2][4] ),
    .A2(net241),
    .B1(net225),
    .B2(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[22][4] ),
    .ZN(_03330_));
 AOI22_X1 _07570_ (.A1(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[6][4] ),
    .A2(net164),
    .B1(net72),
    .B2(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[24][4] ),
    .ZN(_03331_));
 NAND4_X1 _07571_ (.A1(_03328_),
    .A2(_03329_),
    .A3(_03330_),
    .A4(_03331_),
    .ZN(_03332_));
 NOR4_X1 _07572_ (.A1(_03317_),
    .A2(_03322_),
    .A3(_03327_),
    .A4(_03332_),
    .ZN(_03333_));
 OAI21_X1 _07573_ (.A(_01764_),
    .B1(net130),
    .B2(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[0][4] ),
    .ZN(_03334_));
 AOI22_X1 _07574_ (.A1(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[25][4] ),
    .A2(net154),
    .B1(net243),
    .B2(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[2][4] ),
    .ZN(_03335_));
 AOI22_X1 _07575_ (.A1(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[10][4] ),
    .A2(net91),
    .B1(net232),
    .B2(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[11][4] ),
    .ZN(_03336_));
 AOI22_X1 _07576_ (.A1(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[3][4] ),
    .A2(net64),
    .B1(net106),
    .B2(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[15][4] ),
    .ZN(_03337_));
 AOI22_X1 _07577_ (.A1(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[28][4] ),
    .A2(net75),
    .B1(net197),
    .B2(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[19][4] ),
    .ZN(_03338_));
 NAND4_X2 _07578_ (.A1(_03335_),
    .A2(_03336_),
    .A3(_03337_),
    .A4(_03338_),
    .ZN(_03339_));
 AOI22_X1 _07579_ (.A1(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[4][4] ),
    .A2(net125),
    .B1(net257),
    .B2(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[1][4] ),
    .ZN(_03340_));
 AOI22_X1 _07580_ (.A1(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[24][4] ),
    .A2(net72),
    .B1(net86),
    .B2(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[14][4] ),
    .ZN(_03341_));
 AOI22_X1 _07581_ (.A1(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[6][4] ),
    .A2(net161),
    .B1(net247),
    .B2(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[20][4] ),
    .ZN(_03342_));
 AOI21_X1 _07582_ (.A(net113),
    .B1(net220),
    .B2(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[9][4] ),
    .ZN(_03343_));
 NAND4_X2 _07583_ (.A1(_03340_),
    .A2(_03341_),
    .A3(_03342_),
    .A4(_03343_),
    .ZN(_03344_));
 AOI22_X2 _07584_ (.A1(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[29][4] ),
    .A2(net140),
    .B1(net264),
    .B2(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[18][4] ),
    .ZN(_03345_));
 AOI22_X2 _07585_ (.A1(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[17][4] ),
    .A2(net78),
    .B1(net182),
    .B2(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[8][4] ),
    .ZN(_03346_));
 AOI22_X2 _07586_ (.A1(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[5][4] ),
    .A2(net136),
    .B1(net207),
    .B2(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[30][4] ),
    .ZN(_03347_));
 AOI22_X2 _07587_ (.A1(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[23][4] ),
    .A2(net98),
    .B1(net223),
    .B2(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[22][4] ),
    .ZN(_03348_));
 NAND4_X4 _07588_ (.A1(_03345_),
    .A2(_03346_),
    .A3(_03347_),
    .A4(_03348_),
    .ZN(_03349_));
 AOI22_X1 _07589_ (.A1(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[7][4] ),
    .A2(net67),
    .B1(net206),
    .B2(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[13][4] ),
    .ZN(_03350_));
 AOI22_X1 _07590_ (.A1(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[27][4] ),
    .A2(net189),
    .B1(net168),
    .B2(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[26][4] ),
    .ZN(_03351_));
 AOI22_X1 _07591_ (.A1(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[31][4] ),
    .A2(net96),
    .B1(net82),
    .B2(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[21][4] ),
    .ZN(_03352_));
 AOI22_X2 _07592_ (.A1(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[16][4] ),
    .A2(net118),
    .B1(net266),
    .B2(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[12][4] ),
    .ZN(_03353_));
 NAND4_X2 _07593_ (.A1(_03350_),
    .A2(_03351_),
    .A3(_03352_),
    .A4(_03353_),
    .ZN(_03354_));
 NOR4_X4 _07594_ (.A1(_03339_),
    .A2(_03344_),
    .A3(_03349_),
    .A4(_03354_),
    .ZN(_03355_));
 OAI21_X1 _07595_ (.A(_01164_),
    .B1(net130),
    .B2(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[0][4] ),
    .ZN(_03356_));
 OAI22_X1 _07596_ (.A1(_03333_),
    .A2(_03334_),
    .B1(_03355_),
    .B2(_03356_),
    .ZN(_03357_));
 NOR4_X1 _07597_ (.A1(_03221_),
    .A2(_03267_),
    .A3(_03312_),
    .A4(_03357_),
    .ZN(_03358_));
 AOI22_X1 _07598_ (.A1(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[1][4] ),
    .A2(net256),
    .B1(net217),
    .B2(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[9][4] ),
    .ZN(_03359_));
 AOI22_X1 _07599_ (.A1(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[14][4] ),
    .A2(net85),
    .B1(net82),
    .B2(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[21][4] ),
    .ZN(_03360_));
 AOI22_X1 _07600_ (.A1(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[17][4] ),
    .A2(net79),
    .B1(net132),
    .B2(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[5][4] ),
    .ZN(_03361_));
 AOI22_X1 _07601_ (.A1(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[28][4] ),
    .A2(net77),
    .B1(net173),
    .B2(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[26][4] ),
    .ZN(_03362_));
 NAND4_X1 _07602_ (.A1(_03359_),
    .A2(_03360_),
    .A3(_03361_),
    .A4(_03362_),
    .ZN(_03363_));
 AOI22_X1 _07603_ (.A1(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[23][4] ),
    .A2(net100),
    .B1(net95),
    .B2(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[31][4] ),
    .ZN(_03364_));
 AOI22_X1 _07604_ (.A1(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[25][4] ),
    .A2(net153),
    .B1(net74),
    .B2(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[24][4] ),
    .ZN(_03365_));
 AOI22_X1 _07605_ (.A1(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[15][4] ),
    .A2(net107),
    .B1(net204),
    .B2(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[13][4] ),
    .ZN(_03366_));
 AOI21_X1 _07606_ (.A(net113),
    .B1(net64),
    .B2(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[3][4] ),
    .ZN(_03367_));
 NAND4_X1 _07607_ (.A1(_03364_),
    .A2(_03365_),
    .A3(_03366_),
    .A4(_03367_),
    .ZN(_03368_));
 AOI22_X1 _07608_ (.A1(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[8][4] ),
    .A2(net181),
    .B1(net263),
    .B2(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[18][4] ),
    .ZN(_03369_));
 AOI22_X1 _07609_ (.A1(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[6][4] ),
    .A2(net162),
    .B1(net208),
    .B2(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[30][4] ),
    .ZN(_03370_));
 AOI22_X1 _07610_ (.A1(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[29][4] ),
    .A2(net142),
    .B1(net267),
    .B2(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[12][4] ),
    .ZN(_03371_));
 AOI22_X1 _07611_ (.A1(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[7][4] ),
    .A2(net68),
    .B1(net250),
    .B2(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[20][4] ),
    .ZN(_03372_));
 NAND4_X1 _07612_ (.A1(_03369_),
    .A2(_03370_),
    .A3(_03371_),
    .A4(_03372_),
    .ZN(_03373_));
 AOI22_X1 _07613_ (.A1(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[10][4] ),
    .A2(net90),
    .B1(net242),
    .B2(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[2][4] ),
    .ZN(_03374_));
 AOI22_X1 _07614_ (.A1(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[16][4] ),
    .A2(net116),
    .B1(net226),
    .B2(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[22][4] ),
    .ZN(_03375_));
 AOI22_X1 _07615_ (.A1(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[27][4] ),
    .A2(net190),
    .B1(net194),
    .B2(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[19][4] ),
    .ZN(_03376_));
 AOI22_X1 _07616_ (.A1(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[4][4] ),
    .A2(net124),
    .B1(net233),
    .B2(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[11][4] ),
    .ZN(_03377_));
 NAND4_X1 _07617_ (.A1(_03374_),
    .A2(_03375_),
    .A3(_03376_),
    .A4(_03377_),
    .ZN(_03378_));
 OR4_X2 _07618_ (.A1(_03363_),
    .A2(_03368_),
    .A3(_03373_),
    .A4(_03378_),
    .ZN(_03379_));
 OAI21_X1 _07619_ (.A(_03379_),
    .B1(net130),
    .B2(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[0][4] ),
    .ZN(_03380_));
 AOI221_X2 _07620_ (.A(_00907_),
    .B1(_03176_),
    .B2(_03358_),
    .C1(_03380_),
    .C2(_01820_),
    .ZN(\rdata_o_n[4] ));
 AOI22_X1 _07621_ (.A1(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[5][5] ),
    .A2(net131),
    .B1(net123),
    .B2(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[4][5] ),
    .ZN(_03381_));
 AOI22_X1 _07622_ (.A1(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[25][5] ),
    .A2(net152),
    .B1(net90),
    .B2(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[10][5] ),
    .ZN(_03382_));
 AOI22_X1 _07623_ (.A1(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[20][5] ),
    .A2(net250),
    .B1(net204),
    .B2(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[13][5] ),
    .ZN(_03383_));
 AOI22_X1 _07624_ (.A1(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[9][5] ),
    .A2(net217),
    .B1(net193),
    .B2(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[19][5] ),
    .ZN(_03384_));
 NAND4_X1 _07625_ (.A1(_03381_),
    .A2(_03382_),
    .A3(_03383_),
    .A4(_03384_),
    .ZN(_03385_));
 AOI22_X1 _07626_ (.A1(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[3][5] ),
    .A2(net66),
    .B1(net268),
    .B2(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[12][5] ),
    .ZN(_03386_));
 AOI22_X1 _07627_ (.A1(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[8][5] ),
    .A2(net180),
    .B1(net71),
    .B2(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[24][5] ),
    .ZN(_03387_));
 AOI22_X1 _07628_ (.A1(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[26][5] ),
    .A2(net175),
    .B1(net83),
    .B2(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[21][5] ),
    .ZN(_03388_));
 AOI21_X1 _07629_ (.A(net114),
    .B1(net208),
    .B2(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[30][5] ),
    .ZN(_03389_));
 NAND4_X1 _07630_ (.A1(_03386_),
    .A2(_03387_),
    .A3(_03388_),
    .A4(_03389_),
    .ZN(_03390_));
 AOI22_X1 _07631_ (.A1(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[6][5] ),
    .A2(net162),
    .B1(net144),
    .B2(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[29][5] ),
    .ZN(_03391_));
 AOI22_X1 _07632_ (.A1(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[15][5] ),
    .A2(net108),
    .B1(net87),
    .B2(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[14][5] ),
    .ZN(_03392_));
 AOI22_X1 _07633_ (.A1(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[18][5] ),
    .A2(net263),
    .B1(net240),
    .B2(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[2][5] ),
    .ZN(_03393_));
 AOI22_X1 _07634_ (.A1(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[16][5] ),
    .A2(net116),
    .B1(net233),
    .B2(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[11][5] ),
    .ZN(_03394_));
 NAND4_X1 _07635_ (.A1(_03391_),
    .A2(_03392_),
    .A3(_03393_),
    .A4(_03394_),
    .ZN(_03395_));
 AOI22_X1 _07636_ (.A1(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[28][5] ),
    .A2(net76),
    .B1(net254),
    .B2(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[1][5] ),
    .ZN(_03396_));
 AOI22_X1 _07637_ (.A1(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[23][5] ),
    .A2(net100),
    .B1(net68),
    .B2(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[7][5] ),
    .ZN(_03397_));
 AOI22_X1 _07638_ (.A1(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[31][5] ),
    .A2(net93),
    .B1(net222),
    .B2(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[22][5] ),
    .ZN(_03398_));
 AOI22_X2 _07639_ (.A1(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[17][5] ),
    .A2(net79),
    .B1(net188),
    .B2(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[27][5] ),
    .ZN(_03399_));
 NAND4_X2 _07640_ (.A1(_03396_),
    .A2(_03397_),
    .A3(_03398_),
    .A4(_03399_),
    .ZN(_03400_));
 NOR4_X2 _07641_ (.A1(_03385_),
    .A2(_03390_),
    .A3(_03395_),
    .A4(_03400_),
    .ZN(_03401_));
 OAI21_X1 _07642_ (.A(_01401_),
    .B1(net130),
    .B2(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[0][5] ),
    .ZN(_03402_));
 AOI22_X1 _07643_ (.A1(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[23][5] ),
    .A2(net103),
    .B1(net74),
    .B2(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[24][5] ),
    .ZN(_03403_));
 AOI22_X1 _07644_ (.A1(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[1][5] ),
    .A2(net257),
    .B1(net82),
    .B2(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[21][5] ),
    .ZN(_03404_));
 AOI22_X1 _07645_ (.A1(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[25][5] ),
    .A2(net154),
    .B1(net205),
    .B2(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[13][5] ),
    .ZN(_03405_));
 AOI22_X2 _07646_ (.A1(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[29][5] ),
    .A2(net143),
    .B1(net137),
    .B2(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[5][5] ),
    .ZN(_03406_));
 NAND4_X2 _07647_ (.A1(_03403_),
    .A2(_03404_),
    .A3(_03405_),
    .A4(_03406_),
    .ZN(_03407_));
 AOI22_X1 _07648_ (.A1(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[7][5] ),
    .A2(net67),
    .B1(net264),
    .B2(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[18][5] ),
    .ZN(_03408_));
 AOI22_X1 _07649_ (.A1(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[4][5] ),
    .A2(net125),
    .B1(net91),
    .B2(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[10][5] ),
    .ZN(_03409_));
 AOI22_X1 _07650_ (.A1(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[12][5] ),
    .A2(net270),
    .B1(net197),
    .B2(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[19][5] ),
    .ZN(_03410_));
 AOI21_X1 _07651_ (.A(net113),
    .B1(net189),
    .B2(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[27][5] ),
    .ZN(_03411_));
 NAND4_X2 _07652_ (.A1(_03408_),
    .A2(_03409_),
    .A3(_03410_),
    .A4(_03411_),
    .ZN(_03412_));
 AOI22_X1 _07653_ (.A1(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[15][5] ),
    .A2(net106),
    .B1(net184),
    .B2(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[8][5] ),
    .ZN(_03413_));
 AOI22_X1 _07654_ (.A1(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[22][5] ),
    .A2(net225),
    .B1(net210),
    .B2(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[30][5] ),
    .ZN(_03414_));
 AOI22_X1 _07655_ (.A1(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[3][5] ),
    .A2(net64),
    .B1(net169),
    .B2(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[26][5] ),
    .ZN(_03415_));
 AOI22_X1 _07656_ (.A1(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[16][5] ),
    .A2(net118),
    .B1(net75),
    .B2(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[28][5] ),
    .ZN(_03416_));
 NAND4_X1 _07657_ (.A1(_03413_),
    .A2(_03414_),
    .A3(_03415_),
    .A4(_03416_),
    .ZN(_03417_));
 AOI22_X1 _07658_ (.A1(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[17][5] ),
    .A2(net80),
    .B1(net85),
    .B2(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[14][5] ),
    .ZN(_03418_));
 AOI22_X1 _07659_ (.A1(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[31][5] ),
    .A2(net96),
    .B1(net247),
    .B2(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[20][5] ),
    .ZN(_03419_));
 AOI22_X1 _07660_ (.A1(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[2][5] ),
    .A2(net241),
    .B1(net220),
    .B2(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[9][5] ),
    .ZN(_03420_));
 AOI22_X1 _07661_ (.A1(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[6][5] ),
    .A2(net161),
    .B1(net235),
    .B2(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[11][5] ),
    .ZN(_03421_));
 NAND4_X1 _07662_ (.A1(_03418_),
    .A2(_03419_),
    .A3(_03420_),
    .A4(_03421_),
    .ZN(_03422_));
 NOR4_X2 _07663_ (.A1(_03407_),
    .A2(_03412_),
    .A3(_03417_),
    .A4(_03422_),
    .ZN(_03423_));
 OAI21_X1 _07664_ (.A(_01350_),
    .B1(net130),
    .B2(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[0][5] ),
    .ZN(_03424_));
 OAI22_X1 _07665_ (.A1(_03401_),
    .A2(_03402_),
    .B1(_03423_),
    .B2(_03424_),
    .ZN(_03425_));
 INV_X1 _07666_ (.A(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[20][5] ),
    .ZN(_03426_));
 INV_X1 _07667_ (.A(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[11][5] ),
    .ZN(_03427_));
 OAI22_X1 _07668_ (.A1(_03426_),
    .A2(_01691_),
    .B1(_02556_),
    .B2(_03427_),
    .ZN(_03428_));
 AOI221_X2 _07669_ (.A(_03428_),
    .B1(net260),
    .B2(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[1][5] ),
    .C1(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[10][5] ),
    .C2(net90),
    .ZN(_03429_));
 INV_X1 _07670_ (.A(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[25][5] ),
    .ZN(_03430_));
 NAND2_X2 _07671_ (.A1(_00933_),
    .A2(_00939_),
    .ZN(_03431_));
 INV_X1 _07672_ (.A(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[13][5] ),
    .ZN(_03432_));
 OAI22_X2 _07673_ (.A1(_03430_),
    .A2(_01470_),
    .B1(_03431_),
    .B2(_03432_),
    .ZN(_03433_));
 AOI221_X2 _07674_ (.A(_03433_),
    .B1(net66),
    .B2(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[3][5] ),
    .C1(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[30][5] ),
    .C2(net212),
    .ZN(_03434_));
 INV_X1 _07675_ (.A(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[18][5] ),
    .ZN(_03435_));
 NAND4_X2 _07676_ (.A1(net7),
    .A2(_00944_),
    .A3(_00946_),
    .A4(_00926_),
    .ZN(_03436_));
 INV_X1 _07677_ (.A(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[19][5] ),
    .ZN(_03437_));
 OAI22_X1 _07678_ (.A1(_03435_),
    .A2(_02024_),
    .B1(_03436_),
    .B2(_03437_),
    .ZN(_03438_));
 AOI221_X2 _07679_ (.A(_03438_),
    .B1(_01019_),
    .B2(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[17][5] ),
    .C1(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[27][5] ),
    .C2(net192),
    .ZN(_03439_));
 INV_X1 _07680_ (.A(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[15][5] ),
    .ZN(_03440_));
 INV_X1 _07681_ (.A(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[5][5] ),
    .ZN(_03441_));
 OAI22_X1 _07682_ (.A1(_03440_),
    .A2(_01029_),
    .B1(_02238_),
    .B2(_03441_),
    .ZN(_03442_));
 AOI221_X2 _07683_ (.A(_03442_),
    .B1(_01076_),
    .B2(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[7][5] ),
    .C1(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[22][5] ),
    .C2(net226),
    .ZN(_03443_));
 NAND4_X2 _07684_ (.A1(_03429_),
    .A2(_03434_),
    .A3(_03439_),
    .A4(_03443_),
    .ZN(_03444_));
 AOI22_X1 _07685_ (.A1(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[23][5] ),
    .A2(net101),
    .B1(net117),
    .B2(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[16][5] ),
    .ZN(_03445_));
 AOI22_X1 _07686_ (.A1(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[29][5] ),
    .A2(net144),
    .B1(net95),
    .B2(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[31][5] ),
    .ZN(_03446_));
 AND2_X1 _07687_ (.A1(_03445_),
    .A2(_03446_),
    .ZN(_03447_));
 INV_X1 _07688_ (.A(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[2][5] ),
    .ZN(_03448_));
 INV_X1 _07689_ (.A(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[24][5] ),
    .ZN(_03449_));
 OAI33_X1 _07690_ (.A1(_03448_),
    .A2(_00952_),
    .A3(_00962_),
    .B1(_00954_),
    .B2(_00979_),
    .B3(_03449_),
    .ZN(_03450_));
 AOI221_X1 _07691_ (.A(_03450_),
    .B1(net83),
    .B2(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[21][5] ),
    .C1(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[28][5] ),
    .C2(net77),
    .ZN(_03451_));
 AOI22_X1 _07692_ (.A1(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[26][5] ),
    .A2(net173),
    .B1(net162),
    .B2(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[6][5] ),
    .ZN(_03452_));
 AOI22_X1 _07693_ (.A1(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[8][5] ),
    .A2(net178),
    .B1(net217),
    .B2(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[9][5] ),
    .ZN(_03453_));
 AND2_X1 _07694_ (.A1(_03452_),
    .A2(_03453_),
    .ZN(_03454_));
 INV_X1 _07695_ (.A(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[4][5] ),
    .ZN(_03455_));
 OAI21_X1 _07696_ (.A(net130),
    .B1(_00941_),
    .B2(_03455_),
    .ZN(_03456_));
 AOI221_X1 _07697_ (.A(_03456_),
    .B1(net269),
    .B2(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[12][5] ),
    .C1(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[14][5] ),
    .C2(net87),
    .ZN(_03457_));
 NAND4_X1 _07698_ (.A1(_03447_),
    .A2(_03451_),
    .A3(_03454_),
    .A4(_03457_),
    .ZN(_03458_));
 OAI221_X2 _07699_ (.A(_01700_),
    .B1(_03444_),
    .B2(_03458_),
    .C1(net130),
    .C2(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[0][5] ),
    .ZN(_03459_));
 AOI22_X1 _07700_ (.A1(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[21][5] ),
    .A2(net84),
    .B1(net220),
    .B2(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[9][5] ),
    .ZN(_03460_));
 AOI22_X1 _07701_ (.A1(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[26][5] ),
    .A2(net168),
    .B1(net149),
    .B2(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[25][5] ),
    .ZN(_03461_));
 AOI221_X2 _07702_ (.A(_01119_),
    .B1(net160),
    .B2(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[6][5] ),
    .C1(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[15][5] ),
    .C2(net109),
    .ZN(_03462_));
 AOI22_X2 _07703_ (.A1(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[12][5] ),
    .A2(net266),
    .B1(net206),
    .B2(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[13][5] ),
    .ZN(_03463_));
 NAND4_X2 _07704_ (.A1(_03460_),
    .A2(_03461_),
    .A3(_03462_),
    .A4(_03463_),
    .ZN(_03464_));
 AOI22_X1 _07705_ (.A1(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[7][5] ),
    .A2(net67),
    .B1(net91),
    .B2(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[10][5] ),
    .ZN(_03465_));
 AOI22_X1 _07706_ (.A1(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[4][5] ),
    .A2(net128),
    .B1(net87),
    .B2(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[14][5] ),
    .ZN(_03466_));
 AOI22_X1 _07707_ (.A1(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[27][5] ),
    .A2(net191),
    .B1(net264),
    .B2(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[18][5] ),
    .ZN(_03467_));
 AOI22_X2 _07708_ (.A1(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[5][5] ),
    .A2(net136),
    .B1(net207),
    .B2(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[30][5] ),
    .ZN(_03468_));
 NAND4_X2 _07709_ (.A1(_03465_),
    .A2(_03466_),
    .A3(_03467_),
    .A4(_03468_),
    .ZN(_03469_));
 AOI22_X1 _07710_ (.A1(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[16][5] ),
    .A2(net119),
    .B1(net232),
    .B2(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[11][5] ),
    .ZN(_03470_));
 AOI22_X1 _07711_ (.A1(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[17][5] ),
    .A2(net78),
    .B1(net258),
    .B2(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[1][5] ),
    .ZN(_03471_));
 AOI22_X1 _07712_ (.A1(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[2][5] ),
    .A2(net243),
    .B1(net198),
    .B2(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[19][5] ),
    .ZN(_03472_));
 AOI22_X1 _07713_ (.A1(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[28][5] ),
    .A2(net75),
    .B1(net72),
    .B2(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[24][5] ),
    .ZN(_03473_));
 NAND4_X1 _07714_ (.A1(_03470_),
    .A2(_03471_),
    .A3(_03472_),
    .A4(_03473_),
    .ZN(_03474_));
 AOI22_X1 _07715_ (.A1(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[23][5] ),
    .A2(net98),
    .B1(_01149_),
    .B2(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[31][5] ),
    .ZN(_03475_));
 AOI222_X2 _07716_ (.A1(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[29][5] ),
    .A2(net140),
    .B1(net248),
    .B2(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[20][5] ),
    .C1(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[8][5] ),
    .C2(net182),
    .ZN(_03476_));
 AOI22_X1 _07717_ (.A1(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[3][5] ),
    .A2(net65),
    .B1(net223),
    .B2(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[22][5] ),
    .ZN(_03477_));
 NAND3_X1 _07718_ (.A1(_03475_),
    .A2(_03476_),
    .A3(_03477_),
    .ZN(_03478_));
 NOR4_X2 _07719_ (.A1(_03464_),
    .A2(_03469_),
    .A3(_03474_),
    .A4(_03478_),
    .ZN(_03479_));
 OAI21_X1 _07720_ (.A(_00923_),
    .B1(net130),
    .B2(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[0][5] ),
    .ZN(_03480_));
 OAI21_X1 _07721_ (.A(_03459_),
    .B1(_03479_),
    .B2(_03480_),
    .ZN(_03481_));
 AOI22_X1 _07722_ (.A1(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[29][5] ),
    .A2(net141),
    .B1(net89),
    .B2(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[10][5] ),
    .ZN(_03482_));
 AOI22_X1 _07723_ (.A1(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[8][5] ),
    .A2(net185),
    .B1(net203),
    .B2(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[13][5] ),
    .ZN(_03483_));
 AOI22_X1 _07724_ (.A1(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[28][5] ),
    .A2(net76),
    .B1(net148),
    .B2(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[25][5] ),
    .ZN(_03484_));
 AOI22_X1 _07725_ (.A1(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[5][5] ),
    .A2(_01057_),
    .B1(net218),
    .B2(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[9][5] ),
    .ZN(_03485_));
 NAND4_X1 _07726_ (.A1(_03482_),
    .A2(_03483_),
    .A3(_03484_),
    .A4(_03485_),
    .ZN(_03486_));
 AOI22_X1 _07727_ (.A1(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[27][5] ),
    .A2(net187),
    .B1(net127),
    .B2(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[4][5] ),
    .ZN(_03487_));
 AOI22_X1 _07728_ (.A1(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[21][5] ),
    .A2(_00981_),
    .B1(_00996_),
    .B2(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[22][5] ),
    .ZN(_03488_));
 AOI22_X1 _07729_ (.A1(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[24][5] ),
    .A2(net73),
    .B1(net88),
    .B2(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[14][5] ),
    .ZN(_03489_));
 AOI21_X1 _07730_ (.A(net115),
    .B1(net63),
    .B2(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[3][5] ),
    .ZN(_03490_));
 NAND4_X2 _07731_ (.A1(_03487_),
    .A2(_03488_),
    .A3(_03489_),
    .A4(_03490_),
    .ZN(_03491_));
 INV_X1 _07732_ (.A(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[31][5] ),
    .ZN(_03492_));
 INV_X1 _07733_ (.A(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[20][5] ),
    .ZN(_03493_));
 OAI22_X1 _07734_ (.A1(_03492_),
    .A2(_00934_),
    .B1(_01691_),
    .B2(_03493_),
    .ZN(_03494_));
 AOI221_X1 _07735_ (.A(_03494_),
    .B1(net69),
    .B2(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[7][5] ),
    .C1(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[19][5] ),
    .C2(net202),
    .ZN(_03495_));
 AOI22_X1 _07736_ (.A1(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[15][5] ),
    .A2(net111),
    .B1(net165),
    .B2(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[6][5] ),
    .ZN(_03496_));
 AOI22_X1 _07737_ (.A1(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[11][5] ),
    .A2(net230),
    .B1(net216),
    .B2(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[30][5] ),
    .ZN(_03497_));
 AND2_X1 _07738_ (.A1(_03496_),
    .A2(_03497_),
    .ZN(_03498_));
 INV_X1 _07739_ (.A(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[16][5] ),
    .ZN(_03499_));
 INV_X1 _07740_ (.A(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[1][5] ),
    .ZN(_03500_));
 OAI22_X1 _07741_ (.A1(_03499_),
    .A2(_01027_),
    .B1(_01210_),
    .B2(_03500_),
    .ZN(_03501_));
 AOI221_X1 _07742_ (.A(_03501_),
    .B1(net238),
    .B2(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[2][5] ),
    .C1(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[17][5] ),
    .C2(net81),
    .ZN(_03502_));
 AOI22_X1 _07743_ (.A1(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[12][5] ),
    .A2(_00950_),
    .B1(_00964_),
    .B2(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[18][5] ),
    .ZN(_03503_));
 AOI22_X1 _07744_ (.A1(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[23][5] ),
    .A2(net97),
    .B1(net166),
    .B2(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[26][5] ),
    .ZN(_03504_));
 AND2_X1 _07745_ (.A1(_03503_),
    .A2(_03504_),
    .ZN(_03505_));
 NAND4_X1 _07746_ (.A1(_03495_),
    .A2(_03498_),
    .A3(_03502_),
    .A4(_03505_),
    .ZN(_03506_));
 NOR3_X2 _07747_ (.A1(_03486_),
    .A2(_03491_),
    .A3(_03506_),
    .ZN(_03507_));
 OAI21_X1 _07748_ (.A(_01662_),
    .B1(net130),
    .B2(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[0][5] ),
    .ZN(_03508_));
 OAI21_X1 _07749_ (.A(_01406_),
    .B1(_03507_),
    .B2(_03508_),
    .ZN(_03509_));
 AOI22_X1 _07750_ (.A1(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[5][5] ),
    .A2(net137),
    .B1(net124),
    .B2(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[4][5] ),
    .ZN(_03510_));
 AOI22_X1 _07751_ (.A1(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[10][5] ),
    .A2(net91),
    .B1(net241),
    .B2(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[2][5] ),
    .ZN(_03511_));
 AOI22_X1 _07752_ (.A1(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[28][5] ),
    .A2(net75),
    .B1(net82),
    .B2(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[21][5] ),
    .ZN(_03512_));
 AOI22_X1 _07753_ (.A1(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[24][5] ),
    .A2(net74),
    .B1(net195),
    .B2(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[19][5] ),
    .ZN(_03513_));
 NAND4_X1 _07754_ (.A1(_03510_),
    .A2(_03511_),
    .A3(_03512_),
    .A4(_03513_),
    .ZN(_03514_));
 AOI22_X1 _07755_ (.A1(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[25][5] ),
    .A2(net154),
    .B1(net67),
    .B2(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[7][5] ),
    .ZN(_03515_));
 AOI22_X1 _07756_ (.A1(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[29][5] ),
    .A2(net145),
    .B1(net96),
    .B2(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[31][5] ),
    .ZN(_03516_));
 AOI22_X1 _07757_ (.A1(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[8][5] ),
    .A2(net184),
    .B1(net271),
    .B2(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[12][5] ),
    .ZN(_03517_));
 AOI21_X1 _07758_ (.A(net113),
    .B1(net161),
    .B2(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[6][5] ),
    .ZN(_03518_));
 NAND4_X1 _07759_ (.A1(_03515_),
    .A2(_03516_),
    .A3(_03517_),
    .A4(_03518_),
    .ZN(_03519_));
 AOI22_X1 _07760_ (.A1(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[17][5] ),
    .A2(net80),
    .B1(net106),
    .B2(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[15][5] ),
    .ZN(_03520_));
 AOI22_X1 _07761_ (.A1(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[23][5] ),
    .A2(net103),
    .B1(net209),
    .B2(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[30][5] ),
    .ZN(_03521_));
 AOI22_X1 _07762_ (.A1(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[18][5] ),
    .A2(net265),
    .B1(net234),
    .B2(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[11][5] ),
    .ZN(_03522_));
 AOI22_X1 _07763_ (.A1(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[16][5] ),
    .A2(net118),
    .B1(net219),
    .B2(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[9][5] ),
    .ZN(_03523_));
 NAND4_X1 _07764_ (.A1(_03520_),
    .A2(_03521_),
    .A3(_03522_),
    .A4(_03523_),
    .ZN(_03524_));
 AOI22_X1 _07765_ (.A1(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[3][5] ),
    .A2(net64),
    .B1(net224),
    .B2(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[22][5] ),
    .ZN(_03525_));
 AOI22_X1 _07766_ (.A1(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[27][5] ),
    .A2(net189),
    .B1(net169),
    .B2(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[26][5] ),
    .ZN(_03526_));
 AOI22_X1 _07767_ (.A1(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[20][5] ),
    .A2(net247),
    .B1(net205),
    .B2(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[13][5] ),
    .ZN(_03527_));
 AOI22_X1 _07768_ (.A1(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[14][5] ),
    .A2(net85),
    .B1(net259),
    .B2(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[1][5] ),
    .ZN(_03528_));
 NAND4_X1 _07769_ (.A1(_03525_),
    .A2(_03526_),
    .A3(_03527_),
    .A4(_03528_),
    .ZN(_03529_));
 NOR4_X2 _07770_ (.A1(_03514_),
    .A2(_03519_),
    .A3(_03524_),
    .A4(_03529_),
    .ZN(_03530_));
 OAI21_X1 _07771_ (.A(_01169_),
    .B1(net130),
    .B2(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[0][5] ),
    .ZN(_03531_));
 AOI22_X2 _07772_ (.A1(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[7][5] ),
    .A2(net69),
    .B1(net273),
    .B2(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[12][5] ),
    .ZN(_03532_));
 AOI22_X2 _07773_ (.A1(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[15][5] ),
    .A2(net110),
    .B1(net203),
    .B2(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[13][5] ),
    .ZN(_03533_));
 AOI22_X2 _07774_ (.A1(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[22][5] ),
    .A2(net227),
    .B1(net214),
    .B2(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[30][5] ),
    .ZN(_03534_));
 AOI22_X2 _07775_ (.A1(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[10][5] ),
    .A2(_00956_),
    .B1(net199),
    .B2(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[19][5] ),
    .ZN(_03535_));
 NAND4_X4 _07776_ (.A1(_03532_),
    .A2(_03533_),
    .A3(_03534_),
    .A4(_03535_),
    .ZN(_03536_));
 AOI22_X1 _07777_ (.A1(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[3][5] ),
    .A2(_01102_),
    .B1(net229),
    .B2(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[11][5] ),
    .ZN(_03537_));
 AOI22_X1 _07778_ (.A1(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[6][5] ),
    .A2(net157),
    .B1(net133),
    .B2(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[5][5] ),
    .ZN(_03538_));
 MUX2_X1 _07779_ (.A(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[24][5] ),
    .B(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[26][5] ),
    .S(net8),
    .Z(_03539_));
 AOI22_X1 _07780_ (.A1(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[8][5] ),
    .A2(_00939_),
    .B1(_03539_),
    .B2(net1),
    .ZN(_03540_));
 INV_X1 _07781_ (.A(_03540_),
    .ZN(_03541_));
 AOI221_X2 _07782_ (.A(net115),
    .B1(_03541_),
    .B2(_02912_),
    .C1(net102),
    .C2(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[23][5] ),
    .ZN(_03542_));
 NAND3_X1 _07783_ (.A1(_03537_),
    .A2(_03538_),
    .A3(_03542_),
    .ZN(_03543_));
 AOI22_X1 _07784_ (.A1(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[28][5] ),
    .A2(net76),
    .B1(net246),
    .B2(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[20][5] ),
    .ZN(_03544_));
 AOI22_X1 _07785_ (.A1(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[25][5] ),
    .A2(net147),
    .B1(_00964_),
    .B2(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[18][5] ),
    .ZN(_03545_));
 AOI22_X1 _07786_ (.A1(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[4][5] ),
    .A2(net126),
    .B1(net261),
    .B2(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[1][5] ),
    .ZN(_03546_));
 AOI22_X2 _07787_ (.A1(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[17][5] ),
    .A2(net79),
    .B1(net88),
    .B2(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[14][5] ),
    .ZN(_03547_));
 NAND4_X2 _07788_ (.A1(_03544_),
    .A2(_03545_),
    .A3(_03546_),
    .A4(_03547_),
    .ZN(_03548_));
 AOI222_X2 _07789_ (.A1(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[27][5] ),
    .A2(net188),
    .B1(net141),
    .B2(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[29][5] ),
    .C1(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[31][5] ),
    .C2(net93),
    .ZN(_03549_));
 AOI22_X1 _07790_ (.A1(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[21][5] ),
    .A2(net83),
    .B1(net218),
    .B2(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[9][5] ),
    .ZN(_03550_));
 AOI22_X1 _07791_ (.A1(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[16][5] ),
    .A2(net120),
    .B1(net238),
    .B2(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[2][5] ),
    .ZN(_03551_));
 NAND3_X2 _07792_ (.A1(_03549_),
    .A2(_03550_),
    .A3(_03551_),
    .ZN(_03552_));
 NOR4_X4 _07793_ (.A1(_03536_),
    .A2(_03543_),
    .A3(_03548_),
    .A4(_03552_),
    .ZN(_03553_));
 OAI21_X1 _07794_ (.A(_01583_),
    .B1(net130),
    .B2(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[0][5] ),
    .ZN(_03554_));
 OAI22_X1 _07795_ (.A1(_03530_),
    .A2(_03531_),
    .B1(_03553_),
    .B2(_03554_),
    .ZN(_03555_));
 NOR4_X1 _07796_ (.A1(_03425_),
    .A2(_03481_),
    .A3(_03509_),
    .A4(_03555_),
    .ZN(_03556_));
 AOI22_X1 _07797_ (.A1(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[25][5] ),
    .A2(net149),
    .B1(net228),
    .B2(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[22][5] ),
    .ZN(_03557_));
 AOI22_X1 _07798_ (.A1(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[28][5] ),
    .A2(_01032_),
    .B1(net183),
    .B2(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[8][5] ),
    .ZN(_03558_));
 AOI22_X1 _07799_ (.A1(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[24][5] ),
    .A2(net73),
    .B1(net198),
    .B2(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[19][5] ),
    .ZN(_03559_));
 AOI22_X2 _07800_ (.A1(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[6][5] ),
    .A2(net160),
    .B1(net84),
    .B2(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[21][5] ),
    .ZN(_03560_));
 NAND4_X2 _07801_ (.A1(_03557_),
    .A2(_03558_),
    .A3(_03559_),
    .A4(_03560_),
    .ZN(_03561_));
 AOI22_X1 _07802_ (.A1(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[31][5] ),
    .A2(_01149_),
    .B1(net89),
    .B2(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[10][5] ),
    .ZN(_03562_));
 AOI22_X1 _07803_ (.A1(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[18][5] ),
    .A2(net264),
    .B1(_00999_),
    .B2(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[9][5] ),
    .ZN(_03563_));
 AOI22_X1 _07804_ (.A1(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[5][5] ),
    .A2(net139),
    .B1(net206),
    .B2(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[13][5] ),
    .ZN(_03564_));
 NOR2_X1 _07805_ (.A1(net1),
    .A2(net10),
    .ZN(_03565_));
 AND3_X1 _07806_ (.A1(net7),
    .A2(net9),
    .A3(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[7][5] ),
    .ZN(_03566_));
 MUX2_X1 _07807_ (.A(_01641_),
    .B(_03566_),
    .S(net8),
    .Z(_03567_));
 AOI22_X1 _07808_ (.A1(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[27][5] ),
    .A2(_01021_),
    .B1(_03565_),
    .B2(_03567_),
    .ZN(_03568_));
 NAND4_X1 _07809_ (.A1(_03562_),
    .A2(_03563_),
    .A3(_03564_),
    .A4(_03568_),
    .ZN(_03569_));
 AOI22_X1 _07810_ (.A1(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[17][5] ),
    .A2(net78),
    .B1(net65),
    .B2(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[3][5] ),
    .ZN(_03570_));
 AOI22_X1 _07811_ (.A1(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[23][5] ),
    .A2(net98),
    .B1(net253),
    .B2(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[1][5] ),
    .ZN(_03571_));
 AOI22_X1 _07812_ (.A1(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[29][5] ),
    .A2(net146),
    .B1(net128),
    .B2(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[4][5] ),
    .ZN(_03572_));
 AOI22_X1 _07813_ (.A1(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[14][5] ),
    .A2(net87),
    .B1(net237),
    .B2(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[11][5] ),
    .ZN(_03573_));
 NAND4_X1 _07814_ (.A1(_03570_),
    .A2(_03571_),
    .A3(_03572_),
    .A4(_03573_),
    .ZN(_03574_));
 AOI222_X2 _07815_ (.A1(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[12][5] ),
    .A2(net272),
    .B1(net243),
    .B2(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[2][5] ),
    .C1(net211),
    .C2(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[30][5] ),
    .ZN(_03575_));
 AOI22_X1 _07816_ (.A1(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[15][5] ),
    .A2(net109),
    .B1(net171),
    .B2(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[26][5] ),
    .ZN(_03576_));
 AOI22_X1 _07817_ (.A1(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[16][5] ),
    .A2(net119),
    .B1(net252),
    .B2(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[20][5] ),
    .ZN(_03577_));
 NAND3_X1 _07818_ (.A1(_03575_),
    .A2(_03576_),
    .A3(_03577_),
    .ZN(_03578_));
 NOR4_X2 _07819_ (.A1(_03561_),
    .A2(_03569_),
    .A3(_03574_),
    .A4(_03578_),
    .ZN(_03579_));
 OAI21_X2 _07820_ (.A(_01408_),
    .B1(net130),
    .B2(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[0][5] ),
    .ZN(_03580_));
 AOI22_X1 _07821_ (.A1(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[29][5] ),
    .A2(net146),
    .B1(net228),
    .B2(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[22][5] ),
    .ZN(_03581_));
 AOI22_X1 _07822_ (.A1(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[26][5] ),
    .A2(net171),
    .B1(net211),
    .B2(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[30][5] ),
    .ZN(_03582_));
 AND2_X1 _07823_ (.A1(_03581_),
    .A2(_03582_),
    .ZN(_03583_));
 INV_X1 _07824_ (.A(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[31][5] ),
    .ZN(_03584_));
 INV_X1 _07825_ (.A(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[12][5] ),
    .ZN(_03585_));
 OAI22_X1 _07826_ (.A1(_03584_),
    .A2(_00934_),
    .B1(_01426_),
    .B2(_03585_),
    .ZN(_03586_));
 AOI221_X1 _07827_ (.A(_03586_),
    .B1(net128),
    .B2(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[4][5] ),
    .C1(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[28][5] ),
    .C2(_01032_),
    .ZN(_03587_));
 INV_X1 _07828_ (.A(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[2][5] ),
    .ZN(_03588_));
 INV_X1 _07829_ (.A(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[24][5] ),
    .ZN(_03589_));
 OAI33_X1 _07830_ (.A1(_03588_),
    .A2(_00952_),
    .A3(_00962_),
    .B1(_00954_),
    .B2(_00979_),
    .B3(_03589_),
    .ZN(_03590_));
 AOI221_X1 _07831_ (.A(_03590_),
    .B1(net156),
    .B2(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[6][5] ),
    .C1(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[17][5] ),
    .C2(net81),
    .ZN(_03591_));
 AOI22_X1 _07832_ (.A1(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[15][5] ),
    .A2(net112),
    .B1(net201),
    .B2(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[19][5] ),
    .ZN(_03592_));
 AOI21_X1 _07833_ (.A(net115),
    .B1(net121),
    .B2(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[16][5] ),
    .ZN(_03593_));
 AND2_X1 _07834_ (.A1(_03592_),
    .A2(_03593_),
    .ZN(_03594_));
 NAND4_X1 _07835_ (.A1(_03583_),
    .A2(_03587_),
    .A3(_03591_),
    .A4(_03594_),
    .ZN(_03595_));
 AOI22_X1 _07836_ (.A1(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[27][5] ),
    .A2(net186),
    .B1(net176),
    .B2(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[8][5] ),
    .ZN(_03596_));
 AOI22_X1 _07837_ (.A1(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[10][5] ),
    .A2(net89),
    .B1(net264),
    .B2(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[18][5] ),
    .ZN(_03597_));
 AOI22_X1 _07838_ (.A1(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[14][5] ),
    .A2(_00971_),
    .B1(_00999_),
    .B2(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[9][5] ),
    .ZN(_03598_));
 AOI22_X2 _07839_ (.A1(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[1][5] ),
    .A2(net253),
    .B1(net206),
    .B2(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[13][5] ),
    .ZN(_03599_));
 NAND4_X2 _07840_ (.A1(_03596_),
    .A2(_03597_),
    .A3(_03598_),
    .A4(_03599_),
    .ZN(_03600_));
 AOI22_X1 _07841_ (.A1(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[21][5] ),
    .A2(net84),
    .B1(net237),
    .B2(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[11][5] ),
    .ZN(_03601_));
 AOI22_X1 _07842_ (.A1(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[3][5] ),
    .A2(net63),
    .B1(net244),
    .B2(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[20][5] ),
    .ZN(_03602_));
 AOI22_X1 _07843_ (.A1(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[23][5] ),
    .A2(net99),
    .B1(net70),
    .B2(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[7][5] ),
    .ZN(_03603_));
 AOI22_X2 _07844_ (.A1(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[25][5] ),
    .A2(net150),
    .B1(net139),
    .B2(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[5][5] ),
    .ZN(_03604_));
 NAND4_X2 _07845_ (.A1(_03601_),
    .A2(_03602_),
    .A3(_03603_),
    .A4(_03604_),
    .ZN(_03605_));
 NOR3_X2 _07846_ (.A1(_03595_),
    .A2(_03600_),
    .A3(_03605_),
    .ZN(_03606_));
 OAI21_X1 _07847_ (.A(_01731_),
    .B1(_01064_),
    .B2(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[0][5] ),
    .ZN(_03607_));
 OAI22_X4 _07848_ (.A1(_03579_),
    .A2(_03580_),
    .B1(_03606_),
    .B2(_03607_),
    .ZN(_03608_));
 AOI22_X1 _07849_ (.A1(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[16][5] ),
    .A2(net118),
    .B1(net170),
    .B2(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[26][5] ),
    .ZN(_03609_));
 AOI22_X1 _07850_ (.A1(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[29][5] ),
    .A2(net143),
    .B1(net125),
    .B2(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[4][5] ),
    .ZN(_03610_));
 AOI22_X1 _07851_ (.A1(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[24][5] ),
    .A2(net72),
    .B1(net212),
    .B2(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[30][5] ),
    .ZN(_03611_));
 AOI22_X1 _07852_ (.A1(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[14][5] ),
    .A2(net86),
    .B1(net224),
    .B2(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[22][5] ),
    .ZN(_03612_));
 NAND4_X2 _07853_ (.A1(_03609_),
    .A2(_03610_),
    .A3(_03611_),
    .A4(_03612_),
    .ZN(_03613_));
 AOI22_X1 _07854_ (.A1(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[10][5] ),
    .A2(net91),
    .B1(net205),
    .B2(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[13][5] ),
    .ZN(_03614_));
 AOI22_X1 _07855_ (.A1(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[12][5] ),
    .A2(_00950_),
    .B1(_01009_),
    .B2(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[19][5] ),
    .ZN(_03615_));
 AOI22_X1 _07856_ (.A1(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[15][5] ),
    .A2(net108),
    .B1(net83),
    .B2(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[21][5] ),
    .ZN(_03616_));
 AOI21_X1 _07857_ (.A(net114),
    .B1(net265),
    .B2(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[18][5] ),
    .ZN(_03617_));
 NAND4_X1 _07858_ (.A1(_03614_),
    .A2(_03615_),
    .A3(_03616_),
    .A4(_03617_),
    .ZN(_03618_));
 AOI22_X1 _07859_ (.A1(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[5][5] ),
    .A2(net139),
    .B1(net249),
    .B2(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[20][5] ),
    .ZN(_03619_));
 AOI22_X1 _07860_ (.A1(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[25][5] ),
    .A2(_01046_),
    .B1(net221),
    .B2(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[9][5] ),
    .ZN(_03620_));
 AOI22_X1 _07861_ (.A1(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[6][5] ),
    .A2(_01042_),
    .B1(_00975_),
    .B2(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[1][5] ),
    .ZN(_03621_));
 AOI22_X1 _07862_ (.A1(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[7][5] ),
    .A2(_01076_),
    .B1(net95),
    .B2(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[31][5] ),
    .ZN(_03622_));
 NAND4_X1 _07863_ (.A1(_03619_),
    .A2(_03620_),
    .A3(_03621_),
    .A4(_03622_),
    .ZN(_03623_));
 AOI22_X1 _07864_ (.A1(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[17][5] ),
    .A2(net78),
    .B1(net65),
    .B2(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[3][5] ),
    .ZN(_03624_));
 AOI22_X1 _07865_ (.A1(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[28][5] ),
    .A2(net77),
    .B1(_01034_),
    .B2(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[8][5] ),
    .ZN(_03625_));
 AOI22_X1 _07866_ (.A1(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[27][5] ),
    .A2(net192),
    .B1(net242),
    .B2(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[2][5] ),
    .ZN(_03626_));
 AOI22_X1 _07867_ (.A1(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[23][5] ),
    .A2(net104),
    .B1(net236),
    .B2(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[11][5] ),
    .ZN(_03627_));
 NAND4_X1 _07868_ (.A1(_03624_),
    .A2(_03625_),
    .A3(_03626_),
    .A4(_03627_),
    .ZN(_03628_));
 NOR4_X1 _07869_ (.A1(_03613_),
    .A2(_03618_),
    .A3(_03623_),
    .A4(_03628_),
    .ZN(_03629_));
 OAI21_X1 _07870_ (.A(_01764_),
    .B1(net130),
    .B2(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[0][5] ),
    .ZN(_03630_));
 AOI22_X1 _07871_ (.A1(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[23][5] ),
    .A2(net102),
    .B1(net71),
    .B2(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[24][5] ),
    .ZN(_03631_));
 AOI22_X1 _07872_ (.A1(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[28][5] ),
    .A2(net76),
    .B1(net263),
    .B2(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[18][5] ),
    .ZN(_03632_));
 AOI22_X1 _07873_ (.A1(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[21][5] ),
    .A2(net83),
    .B1(net217),
    .B2(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[9][5] ),
    .ZN(_03633_));
 AOI22_X1 _07874_ (.A1(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[31][5] ),
    .A2(net93),
    .B1(net260),
    .B2(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[1][5] ),
    .ZN(_03634_));
 NAND4_X1 _07875_ (.A1(_03631_),
    .A2(_03632_),
    .A3(_03633_),
    .A4(_03634_),
    .ZN(_03635_));
 AOI22_X1 _07876_ (.A1(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[10][5] ),
    .A2(_00956_),
    .B1(net233),
    .B2(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[11][5] ),
    .ZN(_03636_));
 AOI22_X1 _07877_ (.A1(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[15][5] ),
    .A2(net108),
    .B1(net69),
    .B2(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[7][5] ),
    .ZN(_03637_));
 AOI22_X1 _07878_ (.A1(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[20][5] ),
    .A2(net245),
    .B1(net196),
    .B2(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[19][5] ),
    .ZN(_03638_));
 AOI22_X1 _07879_ (.A1(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[17][5] ),
    .A2(net79),
    .B1(net134),
    .B2(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[5][5] ),
    .ZN(_03639_));
 NAND4_X2 _07880_ (.A1(_03636_),
    .A2(_03637_),
    .A3(_03638_),
    .A4(_03639_),
    .ZN(_03640_));
 MUX2_X1 _07881_ (.A(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[12][5] ),
    .B(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[14][5] ),
    .S(net8),
    .Z(_03641_));
 AOI221_X1 _07882_ (.A(net114),
    .B1(net92),
    .B2(_03641_),
    .C1(net213),
    .C2(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[30][5] ),
    .ZN(_03642_));
 AOI22_X1 _07883_ (.A1(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[29][5] ),
    .A2(net144),
    .B1(net240),
    .B2(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[2][5] ),
    .ZN(_03643_));
 AOI22_X1 _07884_ (.A1(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[25][5] ),
    .A2(net148),
    .B1(net126),
    .B2(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[4][5] ),
    .ZN(_03644_));
 AOI22_X1 _07885_ (.A1(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[16][5] ),
    .A2(net120),
    .B1(net178),
    .B2(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[8][5] ),
    .ZN(_03645_));
 NAND4_X1 _07886_ (.A1(_03642_),
    .A2(_03643_),
    .A3(_03644_),
    .A4(_03645_),
    .ZN(_03646_));
 AOI22_X1 _07887_ (.A1(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[6][5] ),
    .A2(net158),
    .B1(net222),
    .B2(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[22][5] ),
    .ZN(_03647_));
 AOI22_X1 _07888_ (.A1(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[27][5] ),
    .A2(net188),
    .B1(net203),
    .B2(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[13][5] ),
    .ZN(_03648_));
 AOI22_X1 _07889_ (.A1(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[3][5] ),
    .A2(net66),
    .B1(net174),
    .B2(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[26][5] ),
    .ZN(_03649_));
 NAND3_X1 _07890_ (.A1(_03647_),
    .A2(_03648_),
    .A3(_03649_),
    .ZN(_03650_));
 NOR4_X2 _07891_ (.A1(_03635_),
    .A2(_03640_),
    .A3(_03646_),
    .A4(_03650_),
    .ZN(_03651_));
 OAI21_X1 _07892_ (.A(_01295_),
    .B1(net130),
    .B2(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[0][5] ),
    .ZN(_03652_));
 OAI22_X1 _07893_ (.A1(_03629_),
    .A2(_03630_),
    .B1(_03651_),
    .B2(_03652_),
    .ZN(_03653_));
 AOI22_X1 _07894_ (.A1(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[25][5] ),
    .A2(net153),
    .B1(net224),
    .B2(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[22][5] ),
    .ZN(_03654_));
 AOI22_X1 _07895_ (.A1(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[28][5] ),
    .A2(net75),
    .B1(net124),
    .B2(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[4][5] ),
    .ZN(_03655_));
 AOI22_X1 _07896_ (.A1(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[6][5] ),
    .A2(net163),
    .B1(net269),
    .B2(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[12][5] ),
    .ZN(_03656_));
 AOI22_X1 _07897_ (.A1(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[23][5] ),
    .A2(net101),
    .B1(net90),
    .B2(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[10][5] ),
    .ZN(_03657_));
 NAND4_X1 _07898_ (.A1(_03654_),
    .A2(_03655_),
    .A3(_03656_),
    .A4(_03657_),
    .ZN(_03658_));
 AOI22_X1 _07899_ (.A1(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[11][5] ),
    .A2(net234),
    .B1(net195),
    .B2(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[19][5] ),
    .ZN(_03659_));
 AOI22_X1 _07900_ (.A1(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[21][5] ),
    .A2(net82),
    .B1(net219),
    .B2(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[9][5] ),
    .ZN(_03660_));
 AOI22_X1 _07901_ (.A1(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[18][5] ),
    .A2(net265),
    .B1(net256),
    .B2(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[1][5] ),
    .ZN(_03661_));
 AOI21_X1 _07902_ (.A(net113),
    .B1(net117),
    .B2(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[16][5] ),
    .ZN(_03662_));
 NAND4_X1 _07903_ (.A1(_03659_),
    .A2(_03660_),
    .A3(_03661_),
    .A4(_03662_),
    .ZN(_03663_));
 AOI22_X1 _07904_ (.A1(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[27][5] ),
    .A2(net190),
    .B1(net179),
    .B2(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[8][5] ),
    .ZN(_03664_));
 AOI22_X1 _07905_ (.A1(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[5][5] ),
    .A2(net132),
    .B1(net68),
    .B2(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[7][5] ),
    .ZN(_03665_));
 AOI22_X1 _07906_ (.A1(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[17][5] ),
    .A2(net80),
    .B1(net64),
    .B2(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[3][5] ),
    .ZN(_03666_));
 AOI22_X2 _07907_ (.A1(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[29][5] ),
    .A2(net142),
    .B1(net209),
    .B2(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[30][5] ),
    .ZN(_03667_));
 NAND4_X2 _07908_ (.A1(_03664_),
    .A2(_03665_),
    .A3(_03666_),
    .A4(_03667_),
    .ZN(_03668_));
 AOI22_X1 _07909_ (.A1(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[26][5] ),
    .A2(net170),
    .B1(net95),
    .B2(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[31][5] ),
    .ZN(_03669_));
 AOI22_X1 _07910_ (.A1(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[15][5] ),
    .A2(net107),
    .B1(net204),
    .B2(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[13][5] ),
    .ZN(_03670_));
 AOI22_X1 _07911_ (.A1(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[20][5] ),
    .A2(net251),
    .B1(net241),
    .B2(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[2][5] ),
    .ZN(_03671_));
 AOI22_X2 _07912_ (.A1(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[24][5] ),
    .A2(net74),
    .B1(net85),
    .B2(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[14][5] ),
    .ZN(_03672_));
 NAND4_X2 _07913_ (.A1(_03669_),
    .A2(_03670_),
    .A3(_03671_),
    .A4(_03672_),
    .ZN(_03673_));
 NOR4_X2 _07914_ (.A1(_03658_),
    .A2(_03663_),
    .A3(_03668_),
    .A4(_03673_),
    .ZN(_03674_));
 OAI21_X1 _07915_ (.A(_01539_),
    .B1(net130),
    .B2(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[0][5] ),
    .ZN(_03675_));
 AOI22_X1 _07916_ (.A1(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[28][5] ),
    .A2(net75),
    .B1(net232),
    .B2(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[11][5] ),
    .ZN(_03676_));
 AOI22_X1 _07917_ (.A1(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[26][5] ),
    .A2(net168),
    .B1(net82),
    .B2(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[21][5] ),
    .ZN(_03677_));
 AOI22_X1 _07918_ (.A1(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[30][5] ),
    .A2(net207),
    .B1(net197),
    .B2(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[19][5] ),
    .ZN(_03678_));
 AOI22_X2 _07919_ (.A1(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[18][5] ),
    .A2(net264),
    .B1(net86),
    .B2(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[14][5] ),
    .ZN(_03679_));
 NAND4_X2 _07920_ (.A1(_03676_),
    .A2(_03677_),
    .A3(_03678_),
    .A4(_03679_),
    .ZN(_03680_));
 AOI22_X1 _07921_ (.A1(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[24][5] ),
    .A2(net72),
    .B1(net206),
    .B2(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[13][5] ),
    .ZN(_03681_));
 AOI22_X1 _07922_ (.A1(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[5][5] ),
    .A2(net138),
    .B1(net67),
    .B2(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[7][5] ),
    .ZN(_03682_));
 AOI22_X2 _07923_ (.A1(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[23][5] ),
    .A2(net103),
    .B1(net257),
    .B2(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[1][5] ),
    .ZN(_03683_));
 AOI21_X1 _07924_ (.A(net113),
    .B1(net220),
    .B2(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[9][5] ),
    .ZN(_03684_));
 NAND4_X2 _07925_ (.A1(_03681_),
    .A2(_03682_),
    .A3(_03683_),
    .A4(_03684_),
    .ZN(_03685_));
 AOI22_X2 _07926_ (.A1(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[17][5] ),
    .A2(net78),
    .B1(net119),
    .B2(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[16][5] ),
    .ZN(_03686_));
 AOI22_X2 _07927_ (.A1(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[6][5] ),
    .A2(net160),
    .B1(net140),
    .B2(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[29][5] ),
    .ZN(_03687_));
 AOI22_X2 _07928_ (.A1(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[10][5] ),
    .A2(net91),
    .B1(net248),
    .B2(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[20][5] ),
    .ZN(_03688_));
 AOI22_X2 _07929_ (.A1(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[8][5] ),
    .A2(net182),
    .B1(net149),
    .B2(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[25][5] ),
    .ZN(_03689_));
 NAND4_X4 _07930_ (.A1(_03686_),
    .A2(_03687_),
    .A3(_03688_),
    .A4(_03689_),
    .ZN(_03690_));
 AOI22_X1 _07931_ (.A1(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[3][5] ),
    .A2(net64),
    .B1(net106),
    .B2(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[15][5] ),
    .ZN(_03691_));
 AOI22_X1 _07932_ (.A1(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[27][5] ),
    .A2(net189),
    .B1(net243),
    .B2(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[2][5] ),
    .ZN(_03692_));
 AOI22_X1 _07933_ (.A1(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[31][5] ),
    .A2(net96),
    .B1(net270),
    .B2(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[12][5] ),
    .ZN(_03693_));
 AOI22_X2 _07934_ (.A1(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[4][5] ),
    .A2(net125),
    .B1(net223),
    .B2(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[22][5] ),
    .ZN(_03694_));
 NAND4_X2 _07935_ (.A1(_03691_),
    .A2(_03692_),
    .A3(_03693_),
    .A4(_03694_),
    .ZN(_03695_));
 NOR4_X4 _07936_ (.A1(_03680_),
    .A2(_03685_),
    .A3(_03690_),
    .A4(_03695_),
    .ZN(_03696_));
 OAI21_X1 _07937_ (.A(_01164_),
    .B1(net130),
    .B2(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[0][5] ),
    .ZN(_03697_));
 OAI22_X2 _07938_ (.A1(_03674_),
    .A2(_03675_),
    .B1(_03696_),
    .B2(_03697_),
    .ZN(_03698_));
 AOI22_X1 _07939_ (.A1(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[16][5] ),
    .A2(net121),
    .B1(_00964_),
    .B2(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[18][5] ),
    .ZN(_03699_));
 AOI22_X1 _07940_ (.A1(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[4][5] ),
    .A2(net129),
    .B1(_00986_),
    .B2(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[20][5] ),
    .ZN(_03700_));
 AND2_X1 _07941_ (.A1(_03699_),
    .A2(_03700_),
    .ZN(_03701_));
 INV_X1 _07942_ (.A(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[23][5] ),
    .ZN(_03702_));
 INV_X1 _07943_ (.A(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[10][5] ),
    .ZN(_03703_));
 OAI33_X1 _07944_ (.A1(_03702_),
    .A2(_00960_),
    .A3(_00980_),
    .B1(_00954_),
    .B2(_00952_),
    .B3(_03703_),
    .ZN(_03704_));
 AOI221_X1 _07945_ (.A(_03704_),
    .B1(net73),
    .B2(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[24][5] ),
    .C1(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[25][5] ),
    .C2(net151),
    .ZN(_03705_));
 INV_X1 _07946_ (.A(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[1][5] ),
    .ZN(_03706_));
 INV_X1 _07947_ (.A(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[13][5] ),
    .ZN(_03707_));
 OAI22_X1 _07948_ (.A1(_03706_),
    .A2(_01210_),
    .B1(_03431_),
    .B2(_03707_),
    .ZN(_03708_));
 AOI221_X1 _07949_ (.A(_03708_),
    .B1(net70),
    .B2(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[7][5] ),
    .C1(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[9][5] ),
    .C2(net221),
    .ZN(_03709_));
 INV_X1 _07950_ (.A(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[27][5] ),
    .ZN(_03710_));
 OAI21_X1 _07951_ (.A(_01064_),
    .B1(_02555_),
    .B2(_03710_),
    .ZN(_03711_));
 AOI221_X1 _07952_ (.A(_03711_),
    .B1(_00996_),
    .B2(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[22][5] ),
    .C1(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[28][5] ),
    .C2(_01032_),
    .ZN(_03712_));
 NAND4_X1 _07953_ (.A1(_03701_),
    .A2(_03705_),
    .A3(_03709_),
    .A4(_03712_),
    .ZN(_03713_));
 AOI22_X1 _07954_ (.A1(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[26][5] ),
    .A2(net172),
    .B1(_01050_),
    .B2(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[29][5] ),
    .ZN(_03714_));
 AOI22_X1 _07955_ (.A1(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[15][5] ),
    .A2(net112),
    .B1(_01149_),
    .B2(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[31][5] ),
    .ZN(_03715_));
 AOI22_X1 _07956_ (.A1(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[8][5] ),
    .A2(net176),
    .B1(_00981_),
    .B2(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[21][5] ),
    .ZN(_03716_));
 AOI22_X2 _07957_ (.A1(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[3][5] ),
    .A2(net63),
    .B1(_00989_),
    .B2(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[2][5] ),
    .ZN(_03717_));
 NAND4_X2 _07958_ (.A1(_03714_),
    .A2(_03715_),
    .A3(_03716_),
    .A4(_03717_),
    .ZN(_03718_));
 AOI22_X1 _07959_ (.A1(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[6][5] ),
    .A2(net159),
    .B1(net135),
    .B2(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[5][5] ),
    .ZN(_03719_));
 AOI22_X1 _07960_ (.A1(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[12][5] ),
    .A2(net274),
    .B1(net88),
    .B2(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[14][5] ),
    .ZN(_03720_));
 AOI22_X1 _07961_ (.A1(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[17][5] ),
    .A2(net81),
    .B1(net200),
    .B2(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[19][5] ),
    .ZN(_03721_));
 AOI22_X1 _07962_ (.A1(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[11][5] ),
    .A2(_00993_),
    .B1(net215),
    .B2(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[30][5] ),
    .ZN(_03722_));
 NAND4_X1 _07963_ (.A1(_03719_),
    .A2(_03720_),
    .A3(_03721_),
    .A4(_03722_),
    .ZN(_03723_));
 NOR3_X2 _07964_ (.A1(_03713_),
    .A2(_03718_),
    .A3(_03723_),
    .ZN(_03724_));
 OAI21_X1 _07965_ (.A(_01502_),
    .B1(net130),
    .B2(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[0][5] ),
    .ZN(_03725_));
 AOI22_X1 _07966_ (.A1(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[6][5] ),
    .A2(net158),
    .B1(net202),
    .B2(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[19][5] ),
    .ZN(_03726_));
 AOI22_X1 _07967_ (.A1(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[25][5] ),
    .A2(net148),
    .B1(net214),
    .B2(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[30][5] ),
    .ZN(_03727_));
 AOI22_X1 _07968_ (.A1(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[2][5] ),
    .A2(net238),
    .B1(net229),
    .B2(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[11][5] ),
    .ZN(_03728_));
 AOI22_X1 _07969_ (.A1(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[5][5] ),
    .A2(net133),
    .B1(net218),
    .B2(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[9][5] ),
    .ZN(_03729_));
 AND4_X1 _07970_ (.A1(_03726_),
    .A2(_03727_),
    .A3(_03728_),
    .A4(_03729_),
    .ZN(_03730_));
 AOI22_X1 _07971_ (.A1(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[1][5] ),
    .A2(net261),
    .B1(net227),
    .B2(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[22][5] ),
    .ZN(_03731_));
 AOI22_X1 _07972_ (.A1(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[28][5] ),
    .A2(net76),
    .B1(net70),
    .B2(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[7][5] ),
    .ZN(_03732_));
 AOI22_X1 _07973_ (.A1(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[8][5] ),
    .A2(net185),
    .B1(net127),
    .B2(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[4][5] ),
    .ZN(_03733_));
 AOI22_X1 _07974_ (.A1(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[23][5] ),
    .A2(net97),
    .B1(_00981_),
    .B2(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[21][5] ),
    .ZN(_03734_));
 AND4_X1 _07975_ (.A1(_03731_),
    .A2(_03732_),
    .A3(_03733_),
    .A4(_03734_),
    .ZN(_03735_));
 INV_X1 _07976_ (.A(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[29][5] ),
    .ZN(_03736_));
 INV_X1 _07977_ (.A(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[31][5] ),
    .ZN(_03737_));
 OAI22_X1 _07978_ (.A1(_03736_),
    .A2(_01425_),
    .B1(_00934_),
    .B2(_03737_),
    .ZN(_03738_));
 AOI221_X1 _07979_ (.A(_03738_),
    .B1(_00956_),
    .B2(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[10][5] ),
    .C1(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[27][5] ),
    .C2(net187),
    .ZN(_03739_));
 MUX2_X1 _07980_ (.A(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[12][5] ),
    .B(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[14][5] ),
    .S(net8),
    .Z(_03740_));
 AOI221_X1 _07981_ (.A(net115),
    .B1(net92),
    .B2(_03740_),
    .C1(net111),
    .C2(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[15][5] ),
    .ZN(_03741_));
 INV_X1 _07982_ (.A(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[20][5] ),
    .ZN(_03742_));
 INV_X1 _07983_ (.A(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[13][5] ),
    .ZN(_03743_));
 OAI22_X1 _07984_ (.A1(_03742_),
    .A2(_01691_),
    .B1(_03431_),
    .B2(_03743_),
    .ZN(_03744_));
 AOI221_X1 _07985_ (.A(_03744_),
    .B1(net81),
    .B2(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[17][5] ),
    .C1(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[18][5] ),
    .C2(_00964_),
    .ZN(_03745_));
 INV_X1 _07986_ (.A(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[16][5] ),
    .ZN(_03746_));
 INV_X1 _07987_ (.A(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[26][5] ),
    .ZN(_03747_));
 OAI22_X1 _07988_ (.A1(_03746_),
    .A2(_01027_),
    .B1(_01203_),
    .B2(_03747_),
    .ZN(_03748_));
 AOI221_X1 _07989_ (.A(_03748_),
    .B1(net63),
    .B2(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[3][5] ),
    .C1(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[24][5] ),
    .C2(_01059_),
    .ZN(_03749_));
 AND4_X1 _07990_ (.A1(_03739_),
    .A2(_03741_),
    .A3(_03745_),
    .A4(_03749_),
    .ZN(_03750_));
 AND3_X1 _07991_ (.A1(_03730_),
    .A2(_03735_),
    .A3(_03750_),
    .ZN(_03751_));
 OAI21_X1 _07992_ (.A(_01623_),
    .B1(net130),
    .B2(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[0][5] ),
    .ZN(_03752_));
 OAI22_X2 _07993_ (.A1(_03724_),
    .A2(_03725_),
    .B1(_03751_),
    .B2(_03752_),
    .ZN(_03753_));
 NOR4_X2 _07994_ (.A1(_03608_),
    .A2(_03653_),
    .A3(_03698_),
    .A4(_03753_),
    .ZN(_03754_));
 AOI22_X1 _07995_ (.A1(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[7][5] ),
    .A2(net68),
    .B1(net217),
    .B2(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[9][5] ),
    .ZN(_03755_));
 AOI22_X1 _07996_ (.A1(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[27][5] ),
    .A2(net190),
    .B1(net267),
    .B2(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[12][5] ),
    .ZN(_03756_));
 AOI22_X1 _07997_ (.A1(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[8][5] ),
    .A2(net179),
    .B1(net153),
    .B2(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[25][5] ),
    .ZN(_03757_));
 AOI22_X1 _07998_ (.A1(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[16][5] ),
    .A2(net116),
    .B1(net173),
    .B2(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[26][5] ),
    .ZN(_03758_));
 NAND4_X1 _07999_ (.A1(_03755_),
    .A2(_03756_),
    .A3(_03757_),
    .A4(_03758_),
    .ZN(_03759_));
 AOI222_X2 _08000_ (.A1(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[15][5] ),
    .A2(net107),
    .B1(net90),
    .B2(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[10][5] ),
    .C1(net142),
    .C2(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[29][5] ),
    .ZN(_03760_));
 AOI22_X1 _08001_ (.A1(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[4][5] ),
    .A2(net123),
    .B1(net250),
    .B2(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[20][5] ),
    .ZN(_03761_));
 AOI22_X1 _08002_ (.A1(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[17][5] ),
    .A2(net79),
    .B1(net71),
    .B2(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[24][5] ),
    .ZN(_03762_));
 NAND3_X1 _08003_ (.A1(_03760_),
    .A2(_03761_),
    .A3(_03762_),
    .ZN(_03763_));
 AOI22_X1 _08004_ (.A1(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[14][5] ),
    .A2(net85),
    .B1(net82),
    .B2(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[21][5] ),
    .ZN(_03764_));
 AOI22_X1 _08005_ (.A1(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[3][5] ),
    .A2(net64),
    .B1(net95),
    .B2(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[31][5] ),
    .ZN(_03765_));
 AOI22_X1 _08006_ (.A1(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[2][5] ),
    .A2(net242),
    .B1(net233),
    .B2(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[11][5] ),
    .ZN(_03766_));
 AOI22_X1 _08007_ (.A1(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[13][5] ),
    .A2(net204),
    .B1(net194),
    .B2(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[19][5] ),
    .ZN(_03767_));
 NAND4_X2 _08008_ (.A1(_03764_),
    .A2(_03765_),
    .A3(_03766_),
    .A4(_03767_),
    .ZN(_03768_));
 AOI22_X1 _08009_ (.A1(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[23][5] ),
    .A2(net100),
    .B1(net162),
    .B2(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[6][5] ),
    .ZN(_03769_));
 AOI22_X1 _08010_ (.A1(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[5][5] ),
    .A2(net131),
    .B1(net263),
    .B2(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[18][5] ),
    .ZN(_03770_));
 AOI22_X1 _08011_ (.A1(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[28][5] ),
    .A2(net76),
    .B1(net226),
    .B2(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[22][5] ),
    .ZN(_03771_));
 AOI22_X2 _08012_ (.A1(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[1][5] ),
    .A2(net255),
    .B1(net208),
    .B2(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[30][5] ),
    .ZN(_03772_));
 NAND4_X2 _08013_ (.A1(_03769_),
    .A2(_03770_),
    .A3(_03771_),
    .A4(_03772_),
    .ZN(_03773_));
 NOR4_X2 _08014_ (.A1(_03759_),
    .A2(_03763_),
    .A3(_03768_),
    .A4(_03773_),
    .ZN(_03774_));
 NAND2_X1 _08015_ (.A1(net130),
    .A2(_03774_),
    .ZN(_03775_));
 OAI21_X1 _08016_ (.A(_03775_),
    .B1(net130),
    .B2(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[0][5] ),
    .ZN(_03776_));
 AOI221_X2 _08017_ (.A(_00907_),
    .B1(_03556_),
    .B2(_03754_),
    .C1(_03776_),
    .C2(_01820_),
    .ZN(\rdata_o_n[5] ));
 INV_X1 _08018_ (.A(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[2][6] ),
    .ZN(_03777_));
 INV_X1 _08019_ (.A(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[22][6] ),
    .ZN(_03778_));
 OAI22_X1 _08020_ (.A1(_03777_),
    .A2(_01211_),
    .B1(_01216_),
    .B2(_03778_),
    .ZN(_03779_));
 AOI221_X1 _08021_ (.A(_03779_),
    .B1(net203),
    .B2(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[13][6] ),
    .C1(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[17][6] ),
    .C2(net81),
    .ZN(_03780_));
 AOI22_X1 _08022_ (.A1(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[25][6] ),
    .A2(net147),
    .B1(net261),
    .B2(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[1][6] ),
    .ZN(_03781_));
 AOI22_X1 _08023_ (.A1(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[27][6] ),
    .A2(net187),
    .B1(net97),
    .B2(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[23][6] ),
    .ZN(_03782_));
 AND2_X1 _08024_ (.A1(_03781_),
    .A2(_03782_),
    .ZN(_03783_));
 AOI22_X1 _08025_ (.A1(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[5][6] ),
    .A2(net133),
    .B1(net230),
    .B2(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[11][6] ),
    .ZN(_03784_));
 AOI22_X1 _08026_ (.A1(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[4][6] ),
    .A2(net127),
    .B1(net214),
    .B2(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[30][6] ),
    .ZN(_03785_));
 AND2_X1 _08027_ (.A1(_03784_),
    .A2(_03785_),
    .ZN(_03786_));
 MUX2_X1 _08028_ (.A(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[24][6] ),
    .B(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[26][6] ),
    .S(net8),
    .Z(_03787_));
 AOI22_X1 _08029_ (.A1(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[8][6] ),
    .A2(_00939_),
    .B1(_03787_),
    .B2(net1),
    .ZN(_03788_));
 INV_X1 _08030_ (.A(_03788_),
    .ZN(_03789_));
 AOI221_X1 _08031_ (.A(net115),
    .B1(_03789_),
    .B2(_02912_),
    .C1(net141),
    .C2(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[29][6] ),
    .ZN(_03790_));
 NAND4_X1 _08032_ (.A1(_03780_),
    .A2(_03783_),
    .A3(_03786_),
    .A4(_03790_),
    .ZN(_03791_));
 AOI22_X1 _08033_ (.A1(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[28][6] ),
    .A2(net76),
    .B1(net273),
    .B2(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[12][6] ),
    .ZN(_03792_));
 AOI22_X1 _08034_ (.A1(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[6][6] ),
    .A2(net157),
    .B1(net88),
    .B2(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[14][6] ),
    .ZN(_03793_));
 AOI22_X1 _08035_ (.A1(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[21][6] ),
    .A2(_00981_),
    .B1(net218),
    .B2(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[9][6] ),
    .ZN(_03794_));
 AOI22_X1 _08036_ (.A1(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[15][6] ),
    .A2(net110),
    .B1(net246),
    .B2(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[20][6] ),
    .ZN(_03795_));
 NAND4_X1 _08037_ (.A1(_03792_),
    .A2(_03793_),
    .A3(_03794_),
    .A4(_03795_),
    .ZN(_03796_));
 AOI222_X2 _08038_ (.A1(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[16][6] ),
    .A2(net122),
    .B1(net69),
    .B2(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[7][6] ),
    .C1(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[3][6] ),
    .C2(_01102_),
    .ZN(_03797_));
 AOI22_X1 _08039_ (.A1(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[31][6] ),
    .A2(net94),
    .B1(net199),
    .B2(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[19][6] ),
    .ZN(_03798_));
 AOI22_X1 _08040_ (.A1(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[10][6] ),
    .A2(net89),
    .B1(_00964_),
    .B2(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[18][6] ),
    .ZN(_03799_));
 NAND3_X1 _08041_ (.A1(_03797_),
    .A2(_03798_),
    .A3(_03799_),
    .ZN(_03800_));
 OR3_X2 _08042_ (.A1(_03791_),
    .A2(_03796_),
    .A3(_03800_),
    .ZN(_03801_));
 OAI21_X1 _08043_ (.A(_01583_),
    .B1(net130),
    .B2(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[0][6] ),
    .ZN(_03802_));
 INV_X1 _08044_ (.A(_03802_),
    .ZN(_03803_));
 AOI22_X1 _08045_ (.A1(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[3][6] ),
    .A2(net64),
    .B1(net225),
    .B2(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[22][6] ),
    .ZN(_03804_));
 AOI22_X1 _08046_ (.A1(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[4][6] ),
    .A2(net125),
    .B1(net243),
    .B2(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[2][6] ),
    .ZN(_03805_));
 AOI22_X1 _08047_ (.A1(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[24][6] ),
    .A2(net72),
    .B1(net197),
    .B2(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[19][6] ),
    .ZN(_03806_));
 AOI22_X1 _08048_ (.A1(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[17][6] ),
    .A2(net80),
    .B1(net184),
    .B2(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[8][6] ),
    .ZN(_03807_));
 NAND4_X1 _08049_ (.A1(_03804_),
    .A2(_03805_),
    .A3(_03806_),
    .A4(_03807_),
    .ZN(_03808_));
 AOI22_X1 _08050_ (.A1(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[12][6] ),
    .A2(net270),
    .B1(net82),
    .B2(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[21][6] ),
    .ZN(_03809_));
 AOI22_X1 _08051_ (.A1(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[26][6] ),
    .A2(net169),
    .B1(net257),
    .B2(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[1][6] ),
    .ZN(_03810_));
 AOI22_X1 _08052_ (.A1(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[7][6] ),
    .A2(net67),
    .B1(net247),
    .B2(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[20][6] ),
    .ZN(_03811_));
 AOI21_X1 _08053_ (.A(net113),
    .B1(net161),
    .B2(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[6][6] ),
    .ZN(_03812_));
 NAND4_X1 _08054_ (.A1(_03809_),
    .A2(_03810_),
    .A3(_03811_),
    .A4(_03812_),
    .ZN(_03813_));
 AOI22_X1 _08055_ (.A1(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[5][6] ),
    .A2(net137),
    .B1(net205),
    .B2(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[13][6] ),
    .ZN(_03814_));
 AOI22_X1 _08056_ (.A1(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[16][6] ),
    .A2(net118),
    .B1(net154),
    .B2(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[25][6] ),
    .ZN(_03815_));
 AOI22_X1 _08057_ (.A1(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[28][6] ),
    .A2(net75),
    .B1(net219),
    .B2(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[9][6] ),
    .ZN(_03816_));
 AOI22_X1 _08058_ (.A1(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[29][6] ),
    .A2(net143),
    .B1(net265),
    .B2(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[18][6] ),
    .ZN(_03817_));
 NAND4_X1 _08059_ (.A1(_03814_),
    .A2(_03815_),
    .A3(_03816_),
    .A4(_03817_),
    .ZN(_03818_));
 AOI22_X1 _08060_ (.A1(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[10][6] ),
    .A2(net91),
    .B1(net85),
    .B2(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[14][6] ),
    .ZN(_03819_));
 AOI22_X1 _08061_ (.A1(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[15][6] ),
    .A2(net106),
    .B1(net210),
    .B2(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[30][6] ),
    .ZN(_03820_));
 AOI22_X1 _08062_ (.A1(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[27][6] ),
    .A2(net189),
    .B1(net103),
    .B2(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[23][6] ),
    .ZN(_03821_));
 AOI22_X1 _08063_ (.A1(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[31][6] ),
    .A2(net96),
    .B1(net235),
    .B2(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[11][6] ),
    .ZN(_03822_));
 NAND4_X1 _08064_ (.A1(_03819_),
    .A2(_03820_),
    .A3(_03821_),
    .A4(_03822_),
    .ZN(_03823_));
 OR4_X2 _08065_ (.A1(_03808_),
    .A2(_03813_),
    .A3(_03818_),
    .A4(_03823_),
    .ZN(_03824_));
 OAI21_X1 _08066_ (.A(_01350_),
    .B1(net130),
    .B2(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[0][6] ),
    .ZN(_03825_));
 INV_X1 _08067_ (.A(_03825_),
    .ZN(_03826_));
 AOI22_X1 _08068_ (.A1(_03801_),
    .A2(_03803_),
    .B1(_03824_),
    .B2(_03826_),
    .ZN(_03827_));
 AOI22_X1 _08069_ (.A1(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[7][6] ),
    .A2(_01076_),
    .B1(net272),
    .B2(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[12][6] ),
    .ZN(_03828_));
 AOI21_X1 _08070_ (.A(_01119_),
    .B1(net198),
    .B2(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[19][6] ),
    .ZN(_03829_));
 AOI22_X1 _08071_ (.A1(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[23][6] ),
    .A2(net98),
    .B1(net264),
    .B2(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[18][6] ),
    .ZN(_03830_));
 AOI22_X1 _08072_ (.A1(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[17][6] ),
    .A2(net78),
    .B1(net192),
    .B2(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[27][6] ),
    .ZN(_03831_));
 AND4_X1 _08073_ (.A1(_03828_),
    .A2(_03829_),
    .A3(_03830_),
    .A4(_03831_),
    .ZN(_03832_));
 AOI22_X1 _08074_ (.A1(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[25][6] ),
    .A2(net150),
    .B1(net146),
    .B2(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[29][6] ),
    .ZN(_03833_));
 AOI22_X1 _08075_ (.A1(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[16][6] ),
    .A2(net119),
    .B1(net87),
    .B2(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[14][6] ),
    .ZN(_03834_));
 AOI22_X1 _08076_ (.A1(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[21][6] ),
    .A2(net84),
    .B1(net211),
    .B2(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[30][6] ),
    .ZN(_03835_));
 AOI22_X1 _08077_ (.A1(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[5][6] ),
    .A2(net139),
    .B1(net225),
    .B2(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[22][6] ),
    .ZN(_03836_));
 AND4_X1 _08078_ (.A1(_03833_),
    .A2(_03834_),
    .A3(_03835_),
    .A4(_03836_),
    .ZN(_03837_));
 AOI22_X1 _08079_ (.A1(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[20][6] ),
    .A2(net252),
    .B1(net206),
    .B2(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[13][6] ),
    .ZN(_03838_));
 AOI22_X1 _08080_ (.A1(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[15][6] ),
    .A2(net109),
    .B1(_00975_),
    .B2(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[1][6] ),
    .ZN(_03839_));
 AND2_X1 _08081_ (.A1(_03838_),
    .A2(_03839_),
    .ZN(_03840_));
 INV_X1 _08082_ (.A(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[6][6] ),
    .ZN(_03841_));
 INV_X1 _08083_ (.A(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[11][6] ),
    .ZN(_03842_));
 OAI22_X1 _08084_ (.A1(_03841_),
    .A2(_01681_),
    .B1(_02556_),
    .B2(_03842_),
    .ZN(_03843_));
 AOI221_X1 _08085_ (.A(_03843_),
    .B1(_00999_),
    .B2(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[9][6] ),
    .C1(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[28][6] ),
    .C2(net77),
    .ZN(_03844_));
 INV_X1 _08086_ (.A(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[8][6] ),
    .ZN(_03845_));
 INV_X1 _08087_ (.A(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[2][6] ),
    .ZN(_03846_));
 OAI22_X1 _08088_ (.A1(_03845_),
    .A2(_03001_),
    .B1(_01211_),
    .B2(_03846_),
    .ZN(_03847_));
 AOI221_X1 _08089_ (.A(_03847_),
    .B1(net128),
    .B2(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[4][6] ),
    .C1(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[10][6] ),
    .C2(net89),
    .ZN(_03848_));
 INV_X1 _08090_ (.A(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[26][6] ),
    .ZN(_03849_));
 INV_X1 _08091_ (.A(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[31][6] ),
    .ZN(_03850_));
 OAI22_X1 _08092_ (.A1(_03849_),
    .A2(_01203_),
    .B1(_00934_),
    .B2(_03850_),
    .ZN(_03851_));
 AOI221_X1 _08093_ (.A(_03851_),
    .B1(net65),
    .B2(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[3][6] ),
    .C1(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[24][6] ),
    .C2(net73),
    .ZN(_03852_));
 AND4_X1 _08094_ (.A1(_03840_),
    .A2(_03844_),
    .A3(_03848_),
    .A4(_03852_),
    .ZN(_03853_));
 NAND3_X2 _08095_ (.A1(_03832_),
    .A2(_03837_),
    .A3(_03853_),
    .ZN(_03854_));
 NOR2_X1 _08096_ (.A1(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[0][6] ),
    .A2(net130),
    .ZN(_03855_));
 NOR3_X2 _08097_ (.A1(_01168_),
    .A2(_01407_),
    .A3(_03855_),
    .ZN(_03856_));
 AOI22_X1 _08098_ (.A1(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[31][6] ),
    .A2(_01149_),
    .B1(_01007_),
    .B2(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[13][6] ),
    .ZN(_03857_));
 AOI22_X1 _08099_ (.A1(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[2][6] ),
    .A2(_00989_),
    .B1(net215),
    .B2(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[30][6] ),
    .ZN(_03858_));
 AOI22_X1 _08100_ (.A1(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[17][6] ),
    .A2(net81),
    .B1(_00971_),
    .B2(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[14][6] ),
    .ZN(_03859_));
 AOI22_X1 _08101_ (.A1(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[26][6] ),
    .A2(net172),
    .B1(_00981_),
    .B2(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[21][6] ),
    .ZN(_03860_));
 NAND4_X1 _08102_ (.A1(_03857_),
    .A2(_03858_),
    .A3(_03859_),
    .A4(_03860_),
    .ZN(_03861_));
 AOI22_X1 _08103_ (.A1(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[23][6] ),
    .A2(net99),
    .B1(net128),
    .B2(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[4][6] ),
    .ZN(_03862_));
 AOI22_X1 _08104_ (.A1(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[25][6] ),
    .A2(net150),
    .B1(net201),
    .B2(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[19][6] ),
    .ZN(_03863_));
 AOI22_X1 _08105_ (.A1(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[10][6] ),
    .A2(net89),
    .B1(net264),
    .B2(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[18][6] ),
    .ZN(_03864_));
 AOI22_X2 _08106_ (.A1(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[15][6] ),
    .A2(net112),
    .B1(net253),
    .B2(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[1][6] ),
    .ZN(_03865_));
 NAND4_X2 _08107_ (.A1(_03862_),
    .A2(_03863_),
    .A3(_03864_),
    .A4(_03865_),
    .ZN(_03866_));
 NOR2_X1 _08108_ (.A1(net1),
    .A2(net9),
    .ZN(_03867_));
 NAND3_X1 _08109_ (.A1(net8),
    .A2(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[11][6] ),
    .A3(_01418_),
    .ZN(_03868_));
 OAI21_X1 _08110_ (.A(_03868_),
    .B1(_00985_),
    .B2(net8),
    .ZN(_03869_));
 AOI222_X2 _08111_ (.A1(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[16][6] ),
    .A2(net121),
    .B1(_03867_),
    .B2(_03869_),
    .C1(net228),
    .C2(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[22][6] ),
    .ZN(_03870_));
 AOI22_X1 _08112_ (.A1(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[8][6] ),
    .A2(net176),
    .B1(net274),
    .B2(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[12][6] ),
    .ZN(_03871_));
 AOI22_X1 _08113_ (.A1(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[29][6] ),
    .A2(_01050_),
    .B1(net73),
    .B2(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[24][6] ),
    .ZN(_03872_));
 NAND3_X1 _08114_ (.A1(_03870_),
    .A2(_03871_),
    .A3(_03872_),
    .ZN(_03873_));
 AOI22_X1 _08115_ (.A1(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[3][6] ),
    .A2(net63),
    .B1(net135),
    .B2(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[5][6] ),
    .ZN(_03874_));
 AOI22_X1 _08116_ (.A1(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[27][6] ),
    .A2(net186),
    .B1(_01032_),
    .B2(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[28][6] ),
    .ZN(_03875_));
 AOI22_X1 _08117_ (.A1(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[6][6] ),
    .A2(net156),
    .B1(net70),
    .B2(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[7][6] ),
    .ZN(_03876_));
 AOI22_X1 _08118_ (.A1(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[20][6] ),
    .A2(net244),
    .B1(_00999_),
    .B2(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[9][6] ),
    .ZN(_03877_));
 NAND4_X2 _08119_ (.A1(_03874_),
    .A2(_03875_),
    .A3(_03876_),
    .A4(_03877_),
    .ZN(_03878_));
 OR4_X4 _08120_ (.A1(_03861_),
    .A2(_03866_),
    .A3(_03873_),
    .A4(_03878_),
    .ZN(_03879_));
 OAI21_X1 _08121_ (.A(_01731_),
    .B1(_01064_),
    .B2(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[0][6] ),
    .ZN(_03880_));
 INV_X1 _08122_ (.A(_03880_),
    .ZN(_03881_));
 AOI22_X4 _08123_ (.A1(_03854_),
    .A2(_03856_),
    .B1(_03879_),
    .B2(_03881_),
    .ZN(_03882_));
 AOI22_X1 _08124_ (.A1(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[8][6] ),
    .A2(net178),
    .B1(net158),
    .B2(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[6][6] ),
    .ZN(_03883_));
 NAND2_X4 _08125_ (.A1(_02036_),
    .A2(_02912_),
    .ZN(_03884_));
 INV_X1 _08126_ (.A(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[10][6] ),
    .ZN(_03885_));
 INV_X1 _08127_ (.A(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[16][6] ),
    .ZN(_03886_));
 OAI221_X1 _08128_ (.A(_03883_),
    .B1(_03884_),
    .B2(_03885_),
    .C1(_03886_),
    .C2(_01027_),
    .ZN(_03887_));
 AOI22_X1 _08129_ (.A1(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[23][6] ),
    .A2(net102),
    .B1(net217),
    .B2(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[9][6] ),
    .ZN(_03888_));
 NAND2_X2 _08130_ (.A1(_02036_),
    .A2(_03010_),
    .ZN(_03889_));
 INV_X1 _08131_ (.A(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[7][6] ),
    .ZN(_03890_));
 INV_X1 _08132_ (.A(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[22][6] ),
    .ZN(_03891_));
 OAI221_X1 _08133_ (.A(_03888_),
    .B1(_03889_),
    .B2(_03890_),
    .C1(_03891_),
    .C2(_01216_),
    .ZN(_03892_));
 AOI22_X1 _08134_ (.A1(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[11][6] ),
    .A2(net229),
    .B1(net203),
    .B2(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[13][6] ),
    .ZN(_03893_));
 AOI22_X1 _08135_ (.A1(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[15][6] ),
    .A2(net110),
    .B1(net133),
    .B2(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[5][6] ),
    .ZN(_03894_));
 MUX2_X1 _08136_ (.A(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[12][6] ),
    .B(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[14][6] ),
    .S(net8),
    .Z(_03895_));
 AOI221_X1 _08137_ (.A(net114),
    .B1(net92),
    .B2(_03895_),
    .C1(net126),
    .C2(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[4][6] ),
    .ZN(_03896_));
 NAND3_X1 _08138_ (.A1(_03893_),
    .A2(_03894_),
    .A3(_03896_),
    .ZN(_03897_));
 NOR3_X1 _08139_ (.A1(_03887_),
    .A2(_03892_),
    .A3(_03897_),
    .ZN(_03898_));
 AOI22_X1 _08140_ (.A1(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[27][6] ),
    .A2(net188),
    .B1(net213),
    .B2(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[30][6] ),
    .ZN(_03899_));
 AOI22_X1 _08141_ (.A1(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[26][6] ),
    .A2(net175),
    .B1(net93),
    .B2(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[31][6] ),
    .ZN(_03900_));
 AOI22_X1 _08142_ (.A1(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[21][6] ),
    .A2(net83),
    .B1(net245),
    .B2(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[20][6] ),
    .ZN(_03901_));
 AOI22_X1 _08143_ (.A1(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[28][6] ),
    .A2(net76),
    .B1(net148),
    .B2(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[25][6] ),
    .ZN(_03902_));
 AND4_X1 _08144_ (.A1(_03899_),
    .A2(_03900_),
    .A3(_03901_),
    .A4(_03902_),
    .ZN(_03903_));
 AOI22_X1 _08145_ (.A1(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[17][6] ),
    .A2(net79),
    .B1(net71),
    .B2(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[24][6] ),
    .ZN(_03904_));
 AOI22_X1 _08146_ (.A1(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[29][6] ),
    .A2(net144),
    .B1(net240),
    .B2(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[2][6] ),
    .ZN(_03905_));
 AOI22_X1 _08147_ (.A1(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[3][6] ),
    .A2(net66),
    .B1(net260),
    .B2(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[1][6] ),
    .ZN(_03906_));
 AOI22_X1 _08148_ (.A1(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[18][6] ),
    .A2(net263),
    .B1(net196),
    .B2(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[19][6] ),
    .ZN(_03907_));
 AND4_X1 _08149_ (.A1(_03904_),
    .A2(_03905_),
    .A3(_03906_),
    .A4(_03907_),
    .ZN(_03908_));
 NAND3_X2 _08150_ (.A1(_03898_),
    .A2(_03903_),
    .A3(_03908_),
    .ZN(_03909_));
 NOR2_X1 _08151_ (.A1(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[0][6] ),
    .A2(net130),
    .ZN(_03910_));
 NOR3_X1 _08152_ (.A1(_00921_),
    .A2(_01168_),
    .A3(_03910_),
    .ZN(_03911_));
 AOI21_X1 _08153_ (.A(_01820_),
    .B1(_03909_),
    .B2(_03911_),
    .ZN(_03912_));
 AOI22_X1 _08154_ (.A1(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[12][6] ),
    .A2(net268),
    .B1(net222),
    .B2(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[22][6] ),
    .ZN(_03913_));
 AOI22_X1 _08155_ (.A1(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[16][6] ),
    .A2(net120),
    .B1(net180),
    .B2(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[8][6] ),
    .ZN(_03914_));
 AOI22_X1 _08156_ (.A1(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[27][6] ),
    .A2(net188),
    .B1(net71),
    .B2(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[24][6] ),
    .ZN(_03915_));
 AOI22_X1 _08157_ (.A1(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[14][6] ),
    .A2(net87),
    .B1(net208),
    .B2(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[30][6] ),
    .ZN(_03916_));
 NAND4_X1 _08158_ (.A1(_03913_),
    .A2(_03914_),
    .A3(_03915_),
    .A4(_03916_),
    .ZN(_03917_));
 AOI22_X1 _08159_ (.A1(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[26][6] ),
    .A2(net175),
    .B1(net240),
    .B2(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[2][6] ),
    .ZN(_03918_));
 AOI22_X1 _08160_ (.A1(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[31][6] ),
    .A2(net93),
    .B1(net255),
    .B2(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[1][6] ),
    .ZN(_03919_));
 AOI22_X1 _08161_ (.A1(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[23][6] ),
    .A2(net100),
    .B1(net76),
    .B2(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[28][6] ),
    .ZN(_03920_));
 AOI21_X1 _08162_ (.A(net114),
    .B1(net193),
    .B2(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[19][6] ),
    .ZN(_03921_));
 NAND4_X1 _08163_ (.A1(_03918_),
    .A2(_03919_),
    .A3(_03920_),
    .A4(_03921_),
    .ZN(_03922_));
 AOI22_X1 _08164_ (.A1(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[3][6] ),
    .A2(net66),
    .B1(net162),
    .B2(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[6][6] ),
    .ZN(_03923_));
 AOI22_X1 _08165_ (.A1(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[25][6] ),
    .A2(net152),
    .B1(net131),
    .B2(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[5][6] ),
    .ZN(_03924_));
 AOI22_X1 _08166_ (.A1(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[17][6] ),
    .A2(net79),
    .B1(net204),
    .B2(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[13][6] ),
    .ZN(_03925_));
 AOI22_X1 _08167_ (.A1(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[4][6] ),
    .A2(net123),
    .B1(net236),
    .B2(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[11][6] ),
    .ZN(_03926_));
 NAND4_X1 _08168_ (.A1(_03923_),
    .A2(_03924_),
    .A3(_03925_),
    .A4(_03926_),
    .ZN(_03927_));
 AOI22_X1 _08169_ (.A1(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[15][6] ),
    .A2(net107),
    .B1(net144),
    .B2(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[29][6] ),
    .ZN(_03928_));
 AOI22_X1 _08170_ (.A1(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[7][6] ),
    .A2(net68),
    .B1(net217),
    .B2(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[9][6] ),
    .ZN(_03929_));
 AOI22_X1 _08171_ (.A1(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[18][6] ),
    .A2(net263),
    .B1(net250),
    .B2(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[20][6] ),
    .ZN(_03930_));
 AOI22_X1 _08172_ (.A1(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[10][6] ),
    .A2(net90),
    .B1(net83),
    .B2(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[21][6] ),
    .ZN(_03931_));
 NAND4_X1 _08173_ (.A1(_03928_),
    .A2(_03929_),
    .A3(_03930_),
    .A4(_03931_),
    .ZN(_03932_));
 OR4_X2 _08174_ (.A1(_03917_),
    .A2(_03922_),
    .A3(_03927_),
    .A4(_03932_),
    .ZN(_03933_));
 OAI21_X1 _08175_ (.A(_01401_),
    .B1(net130),
    .B2(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[0][6] ),
    .ZN(_03934_));
 INV_X1 _08176_ (.A(_03934_),
    .ZN(_03935_));
 AOI22_X1 _08177_ (.A1(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[31][6] ),
    .A2(_01149_),
    .B1(net258),
    .B2(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[1][6] ),
    .ZN(_03936_));
 AOI22_X1 _08178_ (.A1(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[8][6] ),
    .A2(net182),
    .B1(net128),
    .B2(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[4][6] ),
    .ZN(_03937_));
 AOI22_X1 _08179_ (.A1(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[24][6] ),
    .A2(net72),
    .B1(net248),
    .B2(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[20][6] ),
    .ZN(_03938_));
 AOI22_X1 _08180_ (.A1(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[23][6] ),
    .A2(net98),
    .B1(net91),
    .B2(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[10][6] ),
    .ZN(_03939_));
 NAND4_X1 _08181_ (.A1(_03936_),
    .A2(_03937_),
    .A3(_03938_),
    .A4(_03939_),
    .ZN(_03940_));
 AOI22_X1 _08182_ (.A1(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[6][6] ),
    .A2(net160),
    .B1(net264),
    .B2(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[18][6] ),
    .ZN(_03941_));
 AOI22_X1 _08183_ (.A1(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[25][6] ),
    .A2(net149),
    .B1(net223),
    .B2(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[22][6] ),
    .ZN(_03942_));
 AOI22_X1 _08184_ (.A1(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[15][6] ),
    .A2(net109),
    .B1(net207),
    .B2(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[30][6] ),
    .ZN(_03943_));
 AOI21_X1 _08185_ (.A(_01119_),
    .B1(net119),
    .B2(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[16][6] ),
    .ZN(_03944_));
 NAND4_X1 _08186_ (.A1(_03941_),
    .A2(_03942_),
    .A3(_03943_),
    .A4(_03944_),
    .ZN(_03945_));
 AOI22_X1 _08187_ (.A1(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[14][6] ),
    .A2(net86),
    .B1(net243),
    .B2(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[2][6] ),
    .ZN(_03946_));
 AOI22_X1 _08188_ (.A1(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[27][6] ),
    .A2(net191),
    .B1(net266),
    .B2(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[12][6] ),
    .ZN(_03947_));
 AOI22_X1 _08189_ (.A1(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[11][6] ),
    .A2(net232),
    .B1(net206),
    .B2(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[13][6] ),
    .ZN(_03948_));
 AOI22_X1 _08190_ (.A1(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[3][6] ),
    .A2(net65),
    .B1(net168),
    .B2(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[26][6] ),
    .ZN(_03949_));
 NAND4_X1 _08191_ (.A1(_03946_),
    .A2(_03947_),
    .A3(_03948_),
    .A4(_03949_),
    .ZN(_03950_));
 AOI22_X1 _08192_ (.A1(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[5][6] ),
    .A2(net136),
    .B1(net198),
    .B2(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[19][6] ),
    .ZN(_03951_));
 AOI22_X1 _08193_ (.A1(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[17][6] ),
    .A2(net78),
    .B1(net67),
    .B2(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[7][6] ),
    .ZN(_03952_));
 AOI22_X1 _08194_ (.A1(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[28][6] ),
    .A2(net75),
    .B1(net84),
    .B2(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[21][6] ),
    .ZN(_03953_));
 AOI22_X1 _08195_ (.A1(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[29][6] ),
    .A2(net140),
    .B1(net220),
    .B2(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[9][6] ),
    .ZN(_03954_));
 NAND4_X1 _08196_ (.A1(_03951_),
    .A2(_03952_),
    .A3(_03953_),
    .A4(_03954_),
    .ZN(_03955_));
 OR4_X2 _08197_ (.A1(_03940_),
    .A2(_03945_),
    .A3(_03950_),
    .A4(_03955_),
    .ZN(_03956_));
 NOR2_X1 _08198_ (.A1(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[0][6] ),
    .A2(net130),
    .ZN(_03957_));
 NOR3_X1 _08199_ (.A1(_00921_),
    .A2(_00922_),
    .A3(_03957_),
    .ZN(_03958_));
 AOI22_X1 _08200_ (.A1(_03933_),
    .A2(_03935_),
    .B1(_03956_),
    .B2(_03958_),
    .ZN(_03959_));
 AND4_X1 _08201_ (.A1(_03827_),
    .A2(_03882_),
    .A3(_03912_),
    .A4(_03959_),
    .ZN(_03960_));
 AOI22_X1 _08202_ (.A1(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[26][6] ),
    .A2(net175),
    .B1(net148),
    .B2(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[25][6] ),
    .ZN(_03961_));
 AOI22_X1 _08203_ (.A1(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[2][6] ),
    .A2(net242),
    .B1(net203),
    .B2(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[13][6] ),
    .ZN(_03962_));
 AOI22_X1 _08204_ (.A1(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[16][6] ),
    .A2(net120),
    .B1(net134),
    .B2(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[5][6] ),
    .ZN(_03963_));
 AOI22_X1 _08205_ (.A1(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[7][6] ),
    .A2(_01076_),
    .B1(net245),
    .B2(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[20][6] ),
    .ZN(_03964_));
 NAND4_X1 _08206_ (.A1(_03961_),
    .A2(_03962_),
    .A3(_03963_),
    .A4(_03964_),
    .ZN(_03965_));
 AOI22_X1 _08207_ (.A1(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[12][6] ),
    .A2(net269),
    .B1(net226),
    .B2(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[22][6] ),
    .ZN(_03966_));
 AOI22_X1 _08208_ (.A1(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[18][6] ),
    .A2(net263),
    .B1(net196),
    .B2(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[19][6] ),
    .ZN(_03967_));
 AOI22_X1 _08209_ (.A1(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[15][6] ),
    .A2(net108),
    .B1(net87),
    .B2(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[14][6] ),
    .ZN(_03968_));
 AOI21_X1 _08210_ (.A(net114),
    .B1(net218),
    .B2(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[9][6] ),
    .ZN(_03969_));
 NAND4_X1 _08211_ (.A1(_03966_),
    .A2(_03967_),
    .A3(_03968_),
    .A4(_03969_),
    .ZN(_03970_));
 AOI22_X1 _08212_ (.A1(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[3][6] ),
    .A2(net64),
    .B1(net101),
    .B2(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[23][6] ),
    .ZN(_03971_));
 AOI22_X1 _08213_ (.A1(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[17][6] ),
    .A2(net80),
    .B1(net90),
    .B2(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[10][6] ),
    .ZN(_03972_));
 AOI22_X1 _08214_ (.A1(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[8][6] ),
    .A2(net181),
    .B1(net144),
    .B2(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[29][6] ),
    .ZN(_03973_));
 AOI22_X1 _08215_ (.A1(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[6][6] ),
    .A2(net163),
    .B1(net260),
    .B2(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[1][6] ),
    .ZN(_03974_));
 NAND4_X1 _08216_ (.A1(_03971_),
    .A2(_03972_),
    .A3(_03973_),
    .A4(_03974_),
    .ZN(_03975_));
 AOI22_X1 _08217_ (.A1(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[28][6] ),
    .A2(net77),
    .B1(net212),
    .B2(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[30][6] ),
    .ZN(_03976_));
 AOI22_X1 _08218_ (.A1(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[27][6] ),
    .A2(net188),
    .B1(net74),
    .B2(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[24][6] ),
    .ZN(_03977_));
 AOI22_X1 _08219_ (.A1(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[31][6] ),
    .A2(net93),
    .B1(net83),
    .B2(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[21][6] ),
    .ZN(_03978_));
 AOI22_X1 _08220_ (.A1(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[4][6] ),
    .A2(net126),
    .B1(net236),
    .B2(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[11][6] ),
    .ZN(_03979_));
 NAND4_X1 _08221_ (.A1(_03976_),
    .A2(_03977_),
    .A3(_03978_),
    .A4(_03979_),
    .ZN(_03980_));
 NOR4_X1 _08222_ (.A1(_03965_),
    .A2(_03970_),
    .A3(_03975_),
    .A4(_03980_),
    .ZN(_03981_));
 OAI21_X1 _08223_ (.A(_01700_),
    .B1(net130),
    .B2(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[0][6] ),
    .ZN(_03982_));
 OR2_X1 _08224_ (.A1(_03981_),
    .A2(_03982_),
    .ZN(_03983_));
 AOI22_X1 _08225_ (.A1(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[30][6] ),
    .A2(net209),
    .B1(net205),
    .B2(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[13][6] ),
    .ZN(_03984_));
 AOI22_X1 _08226_ (.A1(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[28][6] ),
    .A2(net75),
    .B1(net85),
    .B2(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[14][6] ),
    .ZN(_03985_));
 AOI22_X1 _08227_ (.A1(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[8][6] ),
    .A2(net184),
    .B1(net271),
    .B2(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[12][6] ),
    .ZN(_03986_));
 AOI22_X1 _08228_ (.A1(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[29][6] ),
    .A2(net145),
    .B1(net74),
    .B2(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[24][6] ),
    .ZN(_03987_));
 NAND4_X1 _08229_ (.A1(_03984_),
    .A2(_03985_),
    .A3(_03986_),
    .A4(_03987_),
    .ZN(_03988_));
 AOI22_X1 _08230_ (.A1(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[23][6] ),
    .A2(net103),
    .B1(net259),
    .B2(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[1][6] ),
    .ZN(_03989_));
 AOI22_X1 _08231_ (.A1(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[26][6] ),
    .A2(net169),
    .B1(net195),
    .B2(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[19][6] ),
    .ZN(_03990_));
 AOI22_X1 _08232_ (.A1(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[31][6] ),
    .A2(net96),
    .B1(net241),
    .B2(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[2][6] ),
    .ZN(_03991_));
 AOI21_X1 _08233_ (.A(net113),
    .B1(net124),
    .B2(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[4][6] ),
    .ZN(_03992_));
 NAND4_X1 _08234_ (.A1(_03989_),
    .A2(_03990_),
    .A3(_03991_),
    .A4(_03992_),
    .ZN(_03993_));
 AOI22_X1 _08235_ (.A1(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[16][6] ),
    .A2(net118),
    .B1(net91),
    .B2(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[10][6] ),
    .ZN(_03994_));
 AOI22_X1 _08236_ (.A1(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[21][6] ),
    .A2(net82),
    .B1(net234),
    .B2(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[11][6] ),
    .ZN(_03995_));
 AOI22_X1 _08237_ (.A1(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[6][6] ),
    .A2(net161),
    .B1(net137),
    .B2(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[5][6] ),
    .ZN(_03996_));
 AOI22_X1 _08238_ (.A1(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[27][6] ),
    .A2(net189),
    .B1(net219),
    .B2(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[9][6] ),
    .ZN(_03997_));
 NAND4_X1 _08239_ (.A1(_03994_),
    .A2(_03995_),
    .A3(_03996_),
    .A4(_03997_),
    .ZN(_03998_));
 AOI22_X1 _08240_ (.A1(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[7][6] ),
    .A2(net67),
    .B1(net265),
    .B2(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[18][6] ),
    .ZN(_03999_));
 AOI22_X1 _08241_ (.A1(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[15][6] ),
    .A2(net106),
    .B1(net153),
    .B2(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[25][6] ),
    .ZN(_04000_));
 AOI22_X1 _08242_ (.A1(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[3][6] ),
    .A2(net64),
    .B1(net224),
    .B2(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[22][6] ),
    .ZN(_04001_));
 AOI22_X1 _08243_ (.A1(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[17][6] ),
    .A2(net80),
    .B1(net249),
    .B2(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[20][6] ),
    .ZN(_04002_));
 NAND4_X1 _08244_ (.A1(_03999_),
    .A2(_04000_),
    .A3(_04001_),
    .A4(_04002_),
    .ZN(_04003_));
 OR4_X2 _08245_ (.A1(_03988_),
    .A2(_03993_),
    .A3(_03998_),
    .A4(_04003_),
    .ZN(_04004_));
 OAI21_X1 _08246_ (.A(_01169_),
    .B1(net130),
    .B2(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[0][6] ),
    .ZN(_04005_));
 INV_X1 _08247_ (.A(_04005_),
    .ZN(_04006_));
 AOI22_X1 _08248_ (.A1(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[5][6] ),
    .A2(net135),
    .B1(net215),
    .B2(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[30][6] ),
    .ZN(_04007_));
 AOI22_X1 _08249_ (.A1(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[16][6] ),
    .A2(net121),
    .B1(net176),
    .B2(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[8][6] ),
    .ZN(_04008_));
 AOI22_X1 _08250_ (.A1(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[17][6] ),
    .A2(net81),
    .B1(_00975_),
    .B2(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[1][6] ),
    .ZN(_04009_));
 AOI22_X1 _08251_ (.A1(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[27][6] ),
    .A2(net186),
    .B1(net63),
    .B2(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[3][6] ),
    .ZN(_04010_));
 NAND4_X1 _08252_ (.A1(_04007_),
    .A2(_04008_),
    .A3(_04009_),
    .A4(_04010_),
    .ZN(_04011_));
 AOI22_X1 _08253_ (.A1(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[25][6] ),
    .A2(net151),
    .B1(_01149_),
    .B2(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[31][6] ),
    .ZN(_04012_));
 AOI22_X1 _08254_ (.A1(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[23][6] ),
    .A2(_01144_),
    .B1(_00981_),
    .B2(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[21][6] ),
    .ZN(_04013_));
 AOI22_X1 _08255_ (.A1(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[28][6] ),
    .A2(_01032_),
    .B1(net88),
    .B2(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[14][6] ),
    .ZN(_04014_));
 AOI21_X1 _08256_ (.A(net115),
    .B1(net200),
    .B2(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[19][6] ),
    .ZN(_04015_));
 NAND4_X1 _08257_ (.A1(_04012_),
    .A2(_04013_),
    .A3(_04014_),
    .A4(_04015_),
    .ZN(_04016_));
 AOI22_X1 _08258_ (.A1(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[7][6] ),
    .A2(net70),
    .B1(net274),
    .B2(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[12][6] ),
    .ZN(_04017_));
 AOI22_X1 _08259_ (.A1(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[6][6] ),
    .A2(net156),
    .B1(net228),
    .B2(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[22][6] ),
    .ZN(_04018_));
 AOI22_X1 _08260_ (.A1(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[29][6] ),
    .A2(_01050_),
    .B1(net231),
    .B2(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[11][6] ),
    .ZN(_04019_));
 AOI22_X1 _08261_ (.A1(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[15][6] ),
    .A2(net112),
    .B1(net129),
    .B2(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[4][6] ),
    .ZN(_04020_));
 NAND4_X1 _08262_ (.A1(_04017_),
    .A2(_04018_),
    .A3(_04019_),
    .A4(_04020_),
    .ZN(_04021_));
 AOI22_X1 _08263_ (.A1(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[26][6] ),
    .A2(net167),
    .B1(_01059_),
    .B2(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[24][6] ),
    .ZN(_04022_));
 AOI22_X1 _08264_ (.A1(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[2][6] ),
    .A2(_00989_),
    .B1(net221),
    .B2(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[9][6] ),
    .ZN(_04023_));
 AOI22_X1 _08265_ (.A1(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[10][6] ),
    .A2(net89),
    .B1(_01007_),
    .B2(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[13][6] ),
    .ZN(_04024_));
 AOI22_X1 _08266_ (.A1(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[18][6] ),
    .A2(_00964_),
    .B1(net244),
    .B2(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[20][6] ),
    .ZN(_04025_));
 NAND4_X1 _08267_ (.A1(_04022_),
    .A2(_04023_),
    .A3(_04024_),
    .A4(_04025_),
    .ZN(_04026_));
 OR4_X2 _08268_ (.A1(_04011_),
    .A2(_04016_),
    .A3(_04021_),
    .A4(_04026_),
    .ZN(_04027_));
 OAI21_X1 _08269_ (.A(_01502_),
    .B1(net130),
    .B2(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[0][6] ),
    .ZN(_04028_));
 INV_X1 _08270_ (.A(_04028_),
    .ZN(_04029_));
 AOI22_X1 _08271_ (.A1(_04004_),
    .A2(_04006_),
    .B1(_04027_),
    .B2(_04029_),
    .ZN(_04030_));
 AOI21_X1 _08272_ (.A(net113),
    .B1(net195),
    .B2(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[19][6] ),
    .ZN(_04031_));
 AOI22_X1 _08273_ (.A1(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[3][6] ),
    .A2(net64),
    .B1(net85),
    .B2(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[14][6] ),
    .ZN(_04032_));
 AOI22_X1 _08274_ (.A1(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[16][6] ),
    .A2(net117),
    .B1(net241),
    .B2(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[2][6] ),
    .ZN(_04033_));
 AOI22_X1 _08275_ (.A1(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[8][6] ),
    .A2(net179),
    .B1(net269),
    .B2(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[12][6] ),
    .ZN(_04034_));
 NAND4_X1 _08276_ (.A1(_04031_),
    .A2(_04032_),
    .A3(_04033_),
    .A4(_04034_),
    .ZN(_04035_));
 AOI22_X1 _08277_ (.A1(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[24][6] ),
    .A2(net74),
    .B1(net95),
    .B2(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[31][6] ),
    .ZN(_04036_));
 AOI22_X1 _08278_ (.A1(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[21][6] ),
    .A2(net82),
    .B1(net251),
    .B2(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[20][6] ),
    .ZN(_04037_));
 AOI22_X1 _08279_ (.A1(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[17][6] ),
    .A2(net80),
    .B1(net204),
    .B2(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[13][6] ),
    .ZN(_04038_));
 AOI22_X1 _08280_ (.A1(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[26][6] ),
    .A2(net170),
    .B1(net226),
    .B2(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[22][6] ),
    .ZN(_04039_));
 NAND4_X1 _08281_ (.A1(_04036_),
    .A2(_04037_),
    .A3(_04038_),
    .A4(_04039_),
    .ZN(_04040_));
 OR2_X1 _08282_ (.A1(_04035_),
    .A2(_04040_),
    .ZN(_04041_));
 AOI22_X1 _08283_ (.A1(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[15][6] ),
    .A2(net106),
    .B1(net234),
    .B2(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[11][6] ),
    .ZN(_04042_));
 AOI22_X1 _08284_ (.A1(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[27][6] ),
    .A2(net190),
    .B1(net142),
    .B2(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[29][6] ),
    .ZN(_04043_));
 AOI22_X1 _08285_ (.A1(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[28][6] ),
    .A2(net77),
    .B1(net68),
    .B2(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[7][6] ),
    .ZN(_04044_));
 AOI22_X1 _08286_ (.A1(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[6][6] ),
    .A2(net163),
    .B1(net90),
    .B2(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[10][6] ),
    .ZN(_04045_));
 NAND4_X1 _08287_ (.A1(_04042_),
    .A2(_04043_),
    .A3(_04044_),
    .A4(_04045_),
    .ZN(_04046_));
 AOI22_X1 _08288_ (.A1(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[23][6] ),
    .A2(net101),
    .B1(net153),
    .B2(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[25][6] ),
    .ZN(_04047_));
 AOI22_X1 _08289_ (.A1(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[5][6] ),
    .A2(net132),
    .B1(net124),
    .B2(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[4][6] ),
    .ZN(_04048_));
 AOI22_X1 _08290_ (.A1(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[1][6] ),
    .A2(net256),
    .B1(net219),
    .B2(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[9][6] ),
    .ZN(_04049_));
 AOI22_X1 _08291_ (.A1(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[18][6] ),
    .A2(net265),
    .B1(net209),
    .B2(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[30][6] ),
    .ZN(_04050_));
 NAND4_X1 _08292_ (.A1(_04047_),
    .A2(_04048_),
    .A3(_04049_),
    .A4(_04050_),
    .ZN(_04051_));
 OR2_X1 _08293_ (.A1(_04046_),
    .A2(_04051_),
    .ZN(_04052_));
 OAI221_X1 _08294_ (.A(_01539_),
    .B1(_04041_),
    .B2(_04052_),
    .C1(net130),
    .C2(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[0][6] ),
    .ZN(_04053_));
 OAI21_X1 _08295_ (.A(_01164_),
    .B1(_01064_),
    .B2(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[0][6] ),
    .ZN(_04054_));
 AOI22_X1 _08296_ (.A1(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[8][6] ),
    .A2(net183),
    .B1(net168),
    .B2(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[26][6] ),
    .ZN(_04055_));
 INV_X1 _08297_ (.A(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[16][6] ),
    .ZN(_04056_));
 INV_X1 _08298_ (.A(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[24][6] ),
    .ZN(_04057_));
 NAND2_X2 _08299_ (.A1(_01121_),
    .A2(_02912_),
    .ZN(_04058_));
 OAI221_X1 _08300_ (.A(_04055_),
    .B1(_01027_),
    .B2(_04056_),
    .C1(_04057_),
    .C2(_04058_),
    .ZN(_04059_));
 AOI22_X1 _08301_ (.A1(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[22][6] ),
    .A2(net223),
    .B1(net206),
    .B2(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[13][6] ),
    .ZN(_04060_));
 AOI22_X1 _08302_ (.A1(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[20][6] ),
    .A2(net248),
    .B1(net197),
    .B2(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[19][6] ),
    .ZN(_04061_));
 NAND2_X1 _08303_ (.A1(_04060_),
    .A2(_04061_),
    .ZN(_04062_));
 NAND3_X1 _08304_ (.A1(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[17][6] ),
    .A2(_02035_),
    .A3(_01121_),
    .ZN(_04063_));
 NAND2_X1 _08305_ (.A1(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[1][6] ),
    .A2(net258),
    .ZN(_04064_));
 NAND3_X1 _08306_ (.A1(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[3][6] ),
    .A2(_02035_),
    .A3(_02036_),
    .ZN(_04065_));
 NAND3_X1 _08307_ (.A1(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[14][6] ),
    .A2(_02036_),
    .A3(_03013_),
    .ZN(_04066_));
 NAND4_X1 _08308_ (.A1(_04063_),
    .A2(_04064_),
    .A3(_04065_),
    .A4(_04066_),
    .ZN(_04067_));
 AOI22_X1 _08309_ (.A1(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[12][6] ),
    .A2(net270),
    .B1(net264),
    .B2(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[18][6] ),
    .ZN(_04068_));
 INV_X1 _08310_ (.A(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[10][6] ),
    .ZN(_04069_));
 INV_X1 _08311_ (.A(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[23][6] ),
    .ZN(_04070_));
 OAI221_X1 _08312_ (.A(_04068_),
    .B1(_03884_),
    .B2(_04069_),
    .C1(_04070_),
    .C2(_01417_),
    .ZN(_04071_));
 NOR4_X1 _08313_ (.A1(_04059_),
    .A2(_04062_),
    .A3(_04067_),
    .A4(_04071_),
    .ZN(_04072_));
 AOI22_X1 _08314_ (.A1(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[4][6] ),
    .A2(net125),
    .B1(net232),
    .B2(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[11][6] ),
    .ZN(_04073_));
 AOI22_X1 _08315_ (.A1(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[28][6] ),
    .A2(net75),
    .B1(net67),
    .B2(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[7][6] ),
    .ZN(_04074_));
 INV_X1 _08316_ (.A(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[2][6] ),
    .ZN(_04075_));
 INV_X1 _08317_ (.A(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[9][6] ),
    .ZN(_04076_));
 OAI22_X1 _08318_ (.A1(_04075_),
    .A2(_01211_),
    .B1(_01420_),
    .B2(_04076_),
    .ZN(_04077_));
 AOI221_X1 _08319_ (.A(_04077_),
    .B1(net109),
    .B2(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[15][6] ),
    .C1(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[21][6] ),
    .C2(net82),
    .ZN(_04078_));
 AOI22_X1 _08320_ (.A1(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[27][6] ),
    .A2(net189),
    .B1(net140),
    .B2(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[29][6] ),
    .ZN(_04079_));
 AOI22_X1 _08321_ (.A1(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[25][6] ),
    .A2(net149),
    .B1(net96),
    .B2(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[31][6] ),
    .ZN(_04080_));
 AOI22_X1 _08322_ (.A1(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[6][6] ),
    .A2(net160),
    .B1(net136),
    .B2(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[5][6] ),
    .ZN(_04081_));
 AOI21_X1 _08323_ (.A(_01119_),
    .B1(net207),
    .B2(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[30][6] ),
    .ZN(_04082_));
 AND4_X1 _08324_ (.A1(_04079_),
    .A2(_04080_),
    .A3(_04081_),
    .A4(_04082_),
    .ZN(_04083_));
 AND4_X1 _08325_ (.A1(_04073_),
    .A2(_04074_),
    .A3(_04078_),
    .A4(_04083_),
    .ZN(_04084_));
 AOI21_X2 _08326_ (.A(_04054_),
    .B1(_04072_),
    .B2(_04084_),
    .ZN(_04085_));
 OAI21_X1 _08327_ (.A(_01764_),
    .B1(net130),
    .B2(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[0][6] ),
    .ZN(_04086_));
 AOI22_X1 _08328_ (.A1(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[31][6] ),
    .A2(net94),
    .B1(_00975_),
    .B2(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[1][6] ),
    .ZN(_04087_));
 NAND2_X1 _08329_ (.A1(_02035_),
    .A2(_02036_),
    .ZN(_04088_));
 INV_X1 _08330_ (.A(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[3][6] ),
    .ZN(_04089_));
 INV_X1 _08331_ (.A(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[6][6] ),
    .ZN(_04090_));
 OAI221_X1 _08332_ (.A(_04087_),
    .B1(_04088_),
    .B2(_04089_),
    .C1(_04090_),
    .C2(_01681_),
    .ZN(_04091_));
 AOI22_X1 _08333_ (.A1(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[23][6] ),
    .A2(net104),
    .B1(_01002_),
    .B2(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[30][6] ),
    .ZN(_04092_));
 INV_X1 _08334_ (.A(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[7][6] ),
    .ZN(_04093_));
 INV_X1 _08335_ (.A(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[18][6] ),
    .ZN(_04094_));
 OAI221_X1 _08336_ (.A(_04092_),
    .B1(_03889_),
    .B2(_04093_),
    .C1(_04094_),
    .C2(_02024_),
    .ZN(_04095_));
 AOI22_X1 _08337_ (.A1(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[8][6] ),
    .A2(net181),
    .B1(net236),
    .B2(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[11][6] ),
    .ZN(_04096_));
 INV_X1 _08338_ (.A(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[12][6] ),
    .ZN(_04097_));
 INV_X1 _08339_ (.A(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[28][6] ),
    .ZN(_04098_));
 NAND2_X1 _08340_ (.A1(_01121_),
    .A2(_03013_),
    .ZN(_04099_));
 OAI221_X1 _08341_ (.A(_04096_),
    .B1(_01426_),
    .B2(_04097_),
    .C1(_04098_),
    .C2(_04099_),
    .ZN(_04100_));
 NAND3_X1 _08342_ (.A1(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[21][6] ),
    .A2(_01121_),
    .A3(_03010_),
    .ZN(_04101_));
 NAND2_X1 _08343_ (.A1(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[29][6] ),
    .A2(net145),
    .ZN(_04102_));
 AOI22_X1 _08344_ (.A1(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[4][6] ),
    .A2(_01081_),
    .B1(net241),
    .B2(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[2][6] ),
    .ZN(_04103_));
 NAND3_X1 _08345_ (.A1(_04101_),
    .A2(_04102_),
    .A3(_04103_),
    .ZN(_04104_));
 NOR4_X1 _08346_ (.A1(_04091_),
    .A2(_04095_),
    .A3(_04100_),
    .A4(_04104_),
    .ZN(_04105_));
 INV_X1 _08347_ (.A(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[13][6] ),
    .ZN(_04106_));
 INV_X1 _08348_ (.A(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[24][6] ),
    .ZN(_04107_));
 OAI33_X1 _08349_ (.A1(_04106_),
    .A2(_01005_),
    .A3(_00948_),
    .B1(_00954_),
    .B2(_00979_),
    .B3(_04107_),
    .ZN(_04108_));
 AOI221_X1 _08350_ (.A(_04108_),
    .B1(net87),
    .B2(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[14][6] ),
    .C1(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[20][6] ),
    .C2(net249),
    .ZN(_04109_));
 AOI22_X1 _08351_ (.A1(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[15][6] ),
    .A2(_01123_),
    .B1(net225),
    .B2(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[22][6] ),
    .ZN(_04110_));
 AOI22_X1 _08352_ (.A1(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[27][6] ),
    .A2(net192),
    .B1(net198),
    .B2(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[19][6] ),
    .ZN(_04111_));
 AND2_X1 _08353_ (.A1(_04110_),
    .A2(_04111_),
    .ZN(_04112_));
 AOI22_X1 _08354_ (.A1(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[16][6] ),
    .A2(net119),
    .B1(net155),
    .B2(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[25][6] ),
    .ZN(_04113_));
 AOI22_X1 _08355_ (.A1(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[26][6] ),
    .A2(_01038_),
    .B1(net138),
    .B2(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[5][6] ),
    .ZN(_04114_));
 AND2_X1 _08356_ (.A1(_04113_),
    .A2(_04114_),
    .ZN(_04115_));
 INV_X1 _08357_ (.A(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[10][6] ),
    .ZN(_04116_));
 OAI33_X1 _08358_ (.A1(net9),
    .A2(_00985_),
    .A3(_00948_),
    .B1(_00954_),
    .B2(_00952_),
    .B3(_04116_),
    .ZN(_04117_));
 AOI221_X1 _08359_ (.A(_04117_),
    .B1(net221),
    .B2(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[9][6] ),
    .C1(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[17][6] ),
    .C2(net78),
    .ZN(_04118_));
 AND4_X1 _08360_ (.A1(_04109_),
    .A2(_04112_),
    .A3(_04115_),
    .A4(_04118_),
    .ZN(_04119_));
 AOI21_X1 _08361_ (.A(_04086_),
    .B1(_04105_),
    .B2(_04119_),
    .ZN(_00041_));
 OAI21_X1 _08362_ (.A(_01662_),
    .B1(net130),
    .B2(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[0][6] ),
    .ZN(_00042_));
 AOI22_X1 _08363_ (.A1(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[8][6] ),
    .A2(net185),
    .B1(net245),
    .B2(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[20][6] ),
    .ZN(_00043_));
 AOI22_X1 _08364_ (.A1(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[6][6] ),
    .A2(net158),
    .B1(net221),
    .B2(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[9][6] ),
    .ZN(_00044_));
 NAND2_X1 _08365_ (.A1(_00043_),
    .A2(_00044_),
    .ZN(_00045_));
 AOI22_X1 _08366_ (.A1(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[27][6] ),
    .A2(net187),
    .B1(net141),
    .B2(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[29][6] ),
    .ZN(_00046_));
 INV_X1 _08367_ (.A(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[24][6] ),
    .ZN(_00047_));
 INV_X1 _08368_ (.A(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[28][6] ),
    .ZN(_00048_));
 OAI221_X1 _08369_ (.A(_00046_),
    .B1(_04058_),
    .B2(_00047_),
    .C1(_00048_),
    .C2(_04099_),
    .ZN(_00049_));
 AOI22_X1 _08370_ (.A1(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[5][6] ),
    .A2(_01057_),
    .B1(net94),
    .B2(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[31][6] ),
    .ZN(_00050_));
 INV_X1 _08371_ (.A(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[7][6] ),
    .ZN(_00051_));
 INV_X1 _08372_ (.A(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[10][6] ),
    .ZN(_00052_));
 OAI221_X1 _08373_ (.A(_00050_),
    .B1(_03889_),
    .B2(_00051_),
    .C1(_00052_),
    .C2(_03884_),
    .ZN(_00053_));
 AOI22_X1 _08374_ (.A1(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[15][6] ),
    .A2(net111),
    .B1(net167),
    .B2(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[26][6] ),
    .ZN(_00054_));
 AOI22_X1 _08375_ (.A1(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[4][6] ),
    .A2(net127),
    .B1(_00996_),
    .B2(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[22][6] ),
    .ZN(_00055_));
 NAND2_X1 _08376_ (.A1(_00054_),
    .A2(_00055_),
    .ZN(_00056_));
 NOR4_X1 _08377_ (.A1(_00045_),
    .A2(_00049_),
    .A3(_00053_),
    .A4(_00056_),
    .ZN(_00057_));
 INV_X1 _08378_ (.A(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[17][6] ),
    .ZN(_00058_));
 OAI33_X1 _08379_ (.A1(_00058_),
    .A2(_01015_),
    .A3(_00979_),
    .B1(_00985_),
    .B2(_00948_),
    .B3(net9),
    .ZN(_00059_));
 AOI221_X1 _08380_ (.A(_00059_),
    .B1(net63),
    .B2(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[3][6] ),
    .C1(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[14][6] ),
    .C2(net88),
    .ZN(_00060_));
 AOI22_X1 _08381_ (.A1(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[1][6] ),
    .A2(net262),
    .B1(net216),
    .B2(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[30][6] ),
    .ZN(_00061_));
 AOI22_X1 _08382_ (.A1(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[12][6] ),
    .A2(_00950_),
    .B1(_00964_),
    .B2(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[18][6] ),
    .ZN(_00062_));
 AND2_X1 _08383_ (.A1(_00061_),
    .A2(_00062_),
    .ZN(_00063_));
 INV_X1 _08384_ (.A(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[23][6] ),
    .ZN(_00064_));
 INV_X1 _08385_ (.A(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[11][6] ),
    .ZN(_00065_));
 OAI22_X1 _08386_ (.A1(_00064_),
    .A2(_01417_),
    .B1(_02556_),
    .B2(_00065_),
    .ZN(_00066_));
 AOI221_X1 _08387_ (.A(_00066_),
    .B1(net203),
    .B2(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[13][6] ),
    .C1(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[21][6] ),
    .C2(_00981_),
    .ZN(_00067_));
 AOI22_X1 _08388_ (.A1(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[25][6] ),
    .A2(net151),
    .B1(net239),
    .B2(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[2][6] ),
    .ZN(_00068_));
 AOI22_X1 _08389_ (.A1(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[16][6] ),
    .A2(net122),
    .B1(net202),
    .B2(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[19][6] ),
    .ZN(_00069_));
 AND2_X1 _08390_ (.A1(_00068_),
    .A2(_00069_),
    .ZN(_00070_));
 AND4_X1 _08391_ (.A1(_00060_),
    .A2(_00063_),
    .A3(_00067_),
    .A4(_00070_),
    .ZN(_00071_));
 AOI21_X1 _08392_ (.A(_00042_),
    .B1(_00057_),
    .B2(_00071_),
    .ZN(_00072_));
 OAI21_X1 _08393_ (.A(_01623_),
    .B1(net130),
    .B2(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[0][6] ),
    .ZN(_00073_));
 AOI22_X1 _08394_ (.A1(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[15][6] ),
    .A2(net111),
    .B1(net203),
    .B2(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[13][6] ),
    .ZN(_00074_));
 INV_X1 _08395_ (.A(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[24][6] ),
    .ZN(_00075_));
 INV_X1 _08396_ (.A(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[27][6] ),
    .ZN(_00076_));
 OAI221_X1 _08397_ (.A(_00074_),
    .B1(_04058_),
    .B2(_00075_),
    .C1(_00076_),
    .C2(_02555_),
    .ZN(_00077_));
 AOI22_X1 _08398_ (.A1(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[5][6] ),
    .A2(net133),
    .B1(net126),
    .B2(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[4][6] ),
    .ZN(_00078_));
 INV_X1 _08399_ (.A(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[3][6] ),
    .ZN(_00079_));
 INV_X1 _08400_ (.A(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[11][6] ),
    .ZN(_00080_));
 OAI221_X1 _08401_ (.A(_00078_),
    .B1(_04088_),
    .B2(_00079_),
    .C1(_00080_),
    .C2(_02556_),
    .ZN(_00081_));
 NAND2_X1 _08402_ (.A1(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[30][6] ),
    .A2(net214),
    .ZN(_00082_));
 NAND3_X1 _08403_ (.A1(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[21][6] ),
    .A2(_01121_),
    .A3(_03010_),
    .ZN(_00083_));
 AOI22_X1 _08404_ (.A1(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[25][6] ),
    .A2(net148),
    .B1(net245),
    .B2(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[20][6] ),
    .ZN(_00084_));
 NAND3_X1 _08405_ (.A1(_00082_),
    .A2(_00083_),
    .A3(_00084_),
    .ZN(_00085_));
 NAND3_X1 _08406_ (.A1(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[28][6] ),
    .A2(_01121_),
    .A3(_03013_),
    .ZN(_00086_));
 NAND3_X1 _08407_ (.A1(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[10][6] ),
    .A2(_02036_),
    .A3(_02912_),
    .ZN(_00087_));
 NAND2_X1 _08408_ (.A1(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[9][6] ),
    .A2(net218),
    .ZN(_00088_));
 NAND2_X1 _08409_ (.A1(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[6][6] ),
    .A2(net158),
    .ZN(_00089_));
 NAND4_X1 _08410_ (.A1(_00086_),
    .A2(_00087_),
    .A3(_00088_),
    .A4(_00089_),
    .ZN(_00090_));
 NOR4_X1 _08411_ (.A1(_00077_),
    .A2(_00081_),
    .A3(_00085_),
    .A4(_00090_),
    .ZN(_00091_));
 AOI22_X1 _08412_ (.A1(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[17][6] ),
    .A2(net81),
    .B1(net261),
    .B2(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[1][6] ),
    .ZN(_00092_));
 AOI22_X1 _08413_ (.A1(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[2][6] ),
    .A2(net239),
    .B1(net202),
    .B2(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[19][6] ),
    .ZN(_00093_));
 MUX2_X1 _08414_ (.A(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[12][6] ),
    .B(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[14][6] ),
    .S(net8),
    .Z(_00094_));
 AOI221_X1 _08415_ (.A(net115),
    .B1(net92),
    .B2(_00094_),
    .C1(net69),
    .C2(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[7][6] ),
    .ZN(_00095_));
 AOI22_X1 _08416_ (.A1(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[16][6] ),
    .A2(net122),
    .B1(net227),
    .B2(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[22][6] ),
    .ZN(_00096_));
 AOI22_X1 _08417_ (.A1(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[23][6] ),
    .A2(net97),
    .B1(net177),
    .B2(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[8][6] ),
    .ZN(_00097_));
 AOI22_X1 _08418_ (.A1(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[26][6] ),
    .A2(net166),
    .B1(_00964_),
    .B2(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[18][6] ),
    .ZN(_00098_));
 AOI22_X1 _08419_ (.A1(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[29][6] ),
    .A2(net141),
    .B1(net94),
    .B2(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[31][6] ),
    .ZN(_00099_));
 AND4_X1 _08420_ (.A1(_00096_),
    .A2(_00097_),
    .A3(_00098_),
    .A4(_00099_),
    .ZN(_00100_));
 AND4_X1 _08421_ (.A1(_00092_),
    .A2(_00093_),
    .A3(_00095_),
    .A4(_00100_),
    .ZN(_00101_));
 AOI21_X1 _08422_ (.A(_00073_),
    .B1(_00091_),
    .B2(_00101_),
    .ZN(_00102_));
 NOR4_X1 _08423_ (.A1(_04085_),
    .A2(_00041_),
    .A3(_00072_),
    .A4(_00102_),
    .ZN(_00103_));
 AND4_X1 _08424_ (.A1(_03983_),
    .A2(_04030_),
    .A3(_04053_),
    .A4(_00103_),
    .ZN(_00104_));
 AOI22_X1 _08425_ (.A1(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[7][6] ),
    .A2(net68),
    .B1(net217),
    .B2(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[9][6] ),
    .ZN(_00105_));
 AOI22_X1 _08426_ (.A1(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[27][6] ),
    .A2(net190),
    .B1(net267),
    .B2(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[12][6] ),
    .ZN(_00106_));
 AOI22_X1 _08427_ (.A1(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[8][6] ),
    .A2(net179),
    .B1(net153),
    .B2(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[25][6] ),
    .ZN(_00107_));
 AOI22_X2 _08428_ (.A1(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[16][6] ),
    .A2(net116),
    .B1(net173),
    .B2(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[26][6] ),
    .ZN(_00108_));
 NAND4_X2 _08429_ (.A1(_00105_),
    .A2(_00106_),
    .A3(_00107_),
    .A4(_00108_),
    .ZN(_00109_));
 AOI222_X2 _08430_ (.A1(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[15][6] ),
    .A2(net107),
    .B1(net90),
    .B2(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[10][6] ),
    .C1(net142),
    .C2(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[29][6] ),
    .ZN(_00110_));
 AOI22_X1 _08431_ (.A1(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[4][6] ),
    .A2(net123),
    .B1(net250),
    .B2(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[20][6] ),
    .ZN(_00111_));
 AOI22_X1 _08432_ (.A1(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[17][6] ),
    .A2(net79),
    .B1(net71),
    .B2(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[24][6] ),
    .ZN(_00112_));
 NAND3_X1 _08433_ (.A1(_00110_),
    .A2(_00111_),
    .A3(_00112_),
    .ZN(_00113_));
 AOI22_X1 _08434_ (.A1(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[14][6] ),
    .A2(net85),
    .B1(net82),
    .B2(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[21][6] ),
    .ZN(_00114_));
 AOI22_X1 _08435_ (.A1(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[3][6] ),
    .A2(net64),
    .B1(net95),
    .B2(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[31][6] ),
    .ZN(_00115_));
 AOI22_X1 _08436_ (.A1(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[2][6] ),
    .A2(net242),
    .B1(net233),
    .B2(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[11][6] ),
    .ZN(_00116_));
 AOI22_X1 _08437_ (.A1(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[13][6] ),
    .A2(net204),
    .B1(net194),
    .B2(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[19][6] ),
    .ZN(_00117_));
 NAND4_X1 _08438_ (.A1(_00114_),
    .A2(_00115_),
    .A3(_00116_),
    .A4(_00117_),
    .ZN(_00118_));
 AOI22_X1 _08439_ (.A1(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[23][6] ),
    .A2(net100),
    .B1(net162),
    .B2(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[6][6] ),
    .ZN(_00119_));
 AOI22_X1 _08440_ (.A1(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[5][6] ),
    .A2(net131),
    .B1(net263),
    .B2(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[18][6] ),
    .ZN(_00120_));
 AOI22_X1 _08441_ (.A1(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[28][6] ),
    .A2(net76),
    .B1(net226),
    .B2(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[22][6] ),
    .ZN(_00121_));
 AOI22_X2 _08442_ (.A1(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[1][6] ),
    .A2(net255),
    .B1(net208),
    .B2(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[30][6] ),
    .ZN(_00122_));
 NAND4_X2 _08443_ (.A1(_00119_),
    .A2(_00120_),
    .A3(_00121_),
    .A4(_00122_),
    .ZN(_00123_));
 NOR4_X2 _08444_ (.A1(_00109_),
    .A2(_00113_),
    .A3(_00118_),
    .A4(_00123_),
    .ZN(_00124_));
 NAND2_X1 _08445_ (.A1(net130),
    .A2(_00124_),
    .ZN(_00125_));
 OAI21_X1 _08446_ (.A(_00125_),
    .B1(net130),
    .B2(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[0][6] ),
    .ZN(_00126_));
 AOI221_X2 _08447_ (.A(_00907_),
    .B1(_03960_),
    .B2(_00104_),
    .C1(_00126_),
    .C2(_01820_),
    .ZN(\rdata_o_n[6] ));
 OAI21_X1 _08448_ (.A(_01401_),
    .B1(net130),
    .B2(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[0][7] ),
    .ZN(_00127_));
 AOI22_X1 _08449_ (.A1(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[10][7] ),
    .A2(net90),
    .B1(net208),
    .B2(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[30][7] ),
    .ZN(_00128_));
 AOI22_X1 _08450_ (.A1(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[26][7] ),
    .A2(net175),
    .B1(net93),
    .B2(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[31][7] ),
    .ZN(_00129_));
 AOI22_X1 _08451_ (.A1(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[3][7] ),
    .A2(net66),
    .B1(net240),
    .B2(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[2][7] ),
    .ZN(_00130_));
 AOI22_X1 _08452_ (.A1(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[22][7] ),
    .A2(net222),
    .B1(net193),
    .B2(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[19][7] ),
    .ZN(_00131_));
 NAND4_X1 _08453_ (.A1(_00128_),
    .A2(_00129_),
    .A3(_00130_),
    .A4(_00131_),
    .ZN(_00132_));
 AOI222_X2 _08454_ (.A1(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[23][7] ),
    .A2(net100),
    .B1(net68),
    .B2(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[7][7] ),
    .C1(net233),
    .C2(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[11][7] ),
    .ZN(_00133_));
 AOI22_X1 _08455_ (.A1(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[18][7] ),
    .A2(net263),
    .B1(net250),
    .B2(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[20][7] ),
    .ZN(_00134_));
 AOI22_X1 _08456_ (.A1(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[5][7] ),
    .A2(net131),
    .B1(net255),
    .B2(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[1][7] ),
    .ZN(_00135_));
 NAND3_X1 _08457_ (.A1(_00133_),
    .A2(_00134_),
    .A3(_00135_),
    .ZN(_00136_));
 NOR2_X1 _08458_ (.A1(_00132_),
    .A2(_00136_),
    .ZN(_00137_));
 AOI22_X1 _08459_ (.A1(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[4][7] ),
    .A2(net123),
    .B1(net204),
    .B2(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[13][7] ),
    .ZN(_00138_));
 AOI22_X1 _08460_ (.A1(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[25][7] ),
    .A2(net152),
    .B1(net217),
    .B2(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[9][7] ),
    .ZN(_00139_));
 MUX2_X1 _08461_ (.A(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[12][7] ),
    .B(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[14][7] ),
    .S(net8),
    .Z(_00140_));
 AOI221_X1 _08462_ (.A(net114),
    .B1(net92),
    .B2(_00140_),
    .C1(net144),
    .C2(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[29][7] ),
    .ZN(_00141_));
 NAND3_X1 _08463_ (.A1(_00138_),
    .A2(_00139_),
    .A3(_00141_),
    .ZN(_00142_));
 AOI22_X1 _08464_ (.A1(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[28][7] ),
    .A2(net77),
    .B1(net180),
    .B2(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[8][7] ),
    .ZN(_00143_));
 AOI22_X1 _08465_ (.A1(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[17][7] ),
    .A2(net79),
    .B1(net188),
    .B2(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[27][7] ),
    .ZN(_00144_));
 AOI22_X1 _08466_ (.A1(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[15][7] ),
    .A2(_01418_),
    .B1(_00937_),
    .B2(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[6][7] ),
    .ZN(_00145_));
 NOR3_X2 _08467_ (.A1(_00946_),
    .A2(_00952_),
    .A3(_00145_),
    .ZN(_00146_));
 AOI21_X1 _08468_ (.A(_00146_),
    .B1(net116),
    .B2(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[16][7] ),
    .ZN(_00147_));
 AOI22_X1 _08469_ (.A1(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[24][7] ),
    .A2(net71),
    .B1(net83),
    .B2(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[21][7] ),
    .ZN(_00148_));
 NAND4_X1 _08470_ (.A1(_00143_),
    .A2(_00144_),
    .A3(_00147_),
    .A4(_00148_),
    .ZN(_00149_));
 NOR2_X1 _08471_ (.A1(_00142_),
    .A2(_00149_),
    .ZN(_00150_));
 AOI21_X1 _08472_ (.A(_00127_),
    .B1(_00137_),
    .B2(_00150_),
    .ZN(_00151_));
 AOI22_X1 _08473_ (.A1(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[4][7] ),
    .A2(net124),
    .B1(net82),
    .B2(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[21][7] ),
    .ZN(_00152_));
 AOI22_X1 _08474_ (.A1(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[8][7] ),
    .A2(net184),
    .B1(net249),
    .B2(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[20][7] ),
    .ZN(_00153_));
 AOI22_X1 _08475_ (.A1(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[14][7] ),
    .A2(net85),
    .B1(net205),
    .B2(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[13][7] ),
    .ZN(_00154_));
 AOI22_X1 _08476_ (.A1(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[16][7] ),
    .A2(net118),
    .B1(net265),
    .B2(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[18][7] ),
    .ZN(_00155_));
 NAND4_X1 _08477_ (.A1(_00152_),
    .A2(_00153_),
    .A3(_00154_),
    .A4(_00155_),
    .ZN(_00156_));
 AOI22_X1 _08478_ (.A1(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[1][7] ),
    .A2(net259),
    .B1(net195),
    .B2(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[19][7] ),
    .ZN(_00157_));
 AOI22_X1 _08479_ (.A1(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[17][7] ),
    .A2(net80),
    .B1(net106),
    .B2(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[15][7] ),
    .ZN(_00158_));
 AOI22_X1 _08480_ (.A1(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[28][7] ),
    .A2(net75),
    .B1(net74),
    .B2(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[24][7] ),
    .ZN(_00159_));
 AOI21_X1 _08481_ (.A(net113),
    .B1(net101),
    .B2(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[23][7] ),
    .ZN(_00160_));
 NAND4_X1 _08482_ (.A1(_00157_),
    .A2(_00158_),
    .A3(_00159_),
    .A4(_00160_),
    .ZN(_00161_));
 AOI22_X1 _08483_ (.A1(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[25][7] ),
    .A2(net154),
    .B1(net234),
    .B2(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[11][7] ),
    .ZN(_00162_));
 AOI22_X1 _08484_ (.A1(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[5][7] ),
    .A2(net137),
    .B1(net91),
    .B2(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[10][7] ),
    .ZN(_00163_));
 AOI22_X1 _08485_ (.A1(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[26][7] ),
    .A2(net169),
    .B1(net96),
    .B2(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[31][7] ),
    .ZN(_00164_));
 AOI22_X1 _08486_ (.A1(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[6][7] ),
    .A2(net161),
    .B1(net219),
    .B2(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[9][7] ),
    .ZN(_00165_));
 NAND4_X2 _08487_ (.A1(_00162_),
    .A2(_00163_),
    .A3(_00164_),
    .A4(_00165_),
    .ZN(_00166_));
 AOI22_X1 _08488_ (.A1(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[27][7] ),
    .A2(net190),
    .B1(net241),
    .B2(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[2][7] ),
    .ZN(_00167_));
 AOI22_X1 _08489_ (.A1(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[29][7] ),
    .A2(net145),
    .B1(net210),
    .B2(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[30][7] ),
    .ZN(_00168_));
 AOI22_X1 _08490_ (.A1(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[3][7] ),
    .A2(net64),
    .B1(net271),
    .B2(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[12][7] ),
    .ZN(_00169_));
 AOI22_X1 _08491_ (.A1(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[7][7] ),
    .A2(net67),
    .B1(net224),
    .B2(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[22][7] ),
    .ZN(_00170_));
 NAND4_X1 _08492_ (.A1(_00167_),
    .A2(_00168_),
    .A3(_00169_),
    .A4(_00170_),
    .ZN(_00171_));
 NOR4_X1 _08493_ (.A1(_00156_),
    .A2(_00161_),
    .A3(_00166_),
    .A4(_00171_),
    .ZN(_00172_));
 OAI21_X1 _08494_ (.A(_01169_),
    .B1(net130),
    .B2(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[0][7] ),
    .ZN(_00173_));
 AOI22_X1 _08495_ (.A1(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[28][7] ),
    .A2(net75),
    .B1(net223),
    .B2(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[22][7] ),
    .ZN(_00174_));
 AOI22_X1 _08496_ (.A1(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[27][7] ),
    .A2(net189),
    .B1(net136),
    .B2(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[5][7] ),
    .ZN(_00175_));
 AOI22_X1 _08497_ (.A1(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[3][7] ),
    .A2(net65),
    .B1(net220),
    .B2(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[9][7] ),
    .ZN(_00176_));
 AOI22_X1 _08498_ (.A1(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[31][7] ),
    .A2(net96),
    .B1(net264),
    .B2(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[18][7] ),
    .ZN(_00177_));
 NAND4_X1 _08499_ (.A1(_00174_),
    .A2(_00175_),
    .A3(_00176_),
    .A4(_00177_),
    .ZN(_00178_));
 AOI22_X1 _08500_ (.A1(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[7][7] ),
    .A2(net67),
    .B1(net125),
    .B2(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[4][7] ),
    .ZN(_00179_));
 AOI22_X1 _08501_ (.A1(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[16][7] ),
    .A2(net118),
    .B1(net168),
    .B2(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[26][7] ),
    .ZN(_00180_));
 AOI22_X1 _08502_ (.A1(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[23][7] ),
    .A2(net103),
    .B1(net82),
    .B2(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[21][7] ),
    .ZN(_00181_));
 AOI21_X1 _08503_ (.A(_01119_),
    .B1(net210),
    .B2(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[30][7] ),
    .ZN(_00182_));
 NAND4_X2 _08504_ (.A1(_00179_),
    .A2(_00180_),
    .A3(_00181_),
    .A4(_00182_),
    .ZN(_00183_));
 AOI22_X1 _08505_ (.A1(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[29][7] ),
    .A2(net140),
    .B1(net258),
    .B2(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[1][7] ),
    .ZN(_00184_));
 AOI22_X1 _08506_ (.A1(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[6][7] ),
    .A2(net160),
    .B1(net197),
    .B2(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[19][7] ),
    .ZN(_00185_));
 AOI22_X1 _08507_ (.A1(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[25][7] ),
    .A2(net149),
    .B1(net248),
    .B2(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[20][7] ),
    .ZN(_00186_));
 AOI22_X1 _08508_ (.A1(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[8][7] ),
    .A2(net183),
    .B1(net206),
    .B2(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[13][7] ),
    .ZN(_00187_));
 NAND4_X1 _08509_ (.A1(_00184_),
    .A2(_00185_),
    .A3(_00186_),
    .A4(_00187_),
    .ZN(_00188_));
 AOI22_X1 _08510_ (.A1(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[10][7] ),
    .A2(net91),
    .B1(net232),
    .B2(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[11][7] ),
    .ZN(_00189_));
 AOI22_X1 _08511_ (.A1(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[15][7] ),
    .A2(net109),
    .B1(net72),
    .B2(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[24][7] ),
    .ZN(_00190_));
 AOI22_X1 _08512_ (.A1(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[17][7] ),
    .A2(net78),
    .B1(net243),
    .B2(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[2][7] ),
    .ZN(_00191_));
 AOI22_X1 _08513_ (.A1(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[12][7] ),
    .A2(net266),
    .B1(net86),
    .B2(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[14][7] ),
    .ZN(_00192_));
 NAND4_X1 _08514_ (.A1(_00189_),
    .A2(_00190_),
    .A3(_00191_),
    .A4(_00192_),
    .ZN(_00193_));
 NOR4_X2 _08515_ (.A1(_00178_),
    .A2(_00183_),
    .A3(_00188_),
    .A4(_00193_),
    .ZN(_00194_));
 OAI21_X1 _08516_ (.A(_01164_),
    .B1(net130),
    .B2(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[0][7] ),
    .ZN(_00195_));
 OAI22_X1 _08517_ (.A1(_00172_),
    .A2(_00173_),
    .B1(_00194_),
    .B2(_00195_),
    .ZN(_00196_));
 AOI22_X1 _08518_ (.A1(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[16][7] ),
    .A2(net122),
    .B1(net166),
    .B2(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[26][7] ),
    .ZN(_00197_));
 AOI22_X1 _08519_ (.A1(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[6][7] ),
    .A2(net165),
    .B1(_01059_),
    .B2(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[24][7] ),
    .ZN(_00198_));
 AOI22_X1 _08520_ (.A1(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[25][7] ),
    .A2(net147),
    .B1(net141),
    .B2(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[29][7] ),
    .ZN(_00199_));
 AOI22_X1 _08521_ (.A1(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[9][7] ),
    .A2(net218),
    .B1(net216),
    .B2(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[30][7] ),
    .ZN(_00200_));
 NAND4_X1 _08522_ (.A1(_00197_),
    .A2(_00198_),
    .A3(_00199_),
    .A4(_00200_),
    .ZN(_00201_));
 AOI22_X1 _08523_ (.A1(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[27][7] ),
    .A2(net187),
    .B1(net185),
    .B2(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[8][7] ),
    .ZN(_00202_));
 AOI22_X1 _08524_ (.A1(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[31][7] ),
    .A2(net94),
    .B1(net89),
    .B2(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[10][7] ),
    .ZN(_00203_));
 MUX2_X1 _08525_ (.A(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[5][7] ),
    .B(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[21][7] ),
    .S(net1),
    .Z(_00204_));
 AOI221_X1 _08526_ (.A(net115),
    .B1(_01597_),
    .B2(_00204_),
    .C1(net273),
    .C2(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[12][7] ),
    .ZN(_00205_));
 NAND3_X1 _08527_ (.A1(_00202_),
    .A2(_00203_),
    .A3(_00205_),
    .ZN(_00206_));
 AOI22_X1 _08528_ (.A1(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[7][7] ),
    .A2(net70),
    .B1(net239),
    .B2(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[2][7] ),
    .ZN(_00207_));
 AOI22_X1 _08529_ (.A1(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[23][7] ),
    .A2(net97),
    .B1(net127),
    .B2(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[4][7] ),
    .ZN(_00208_));
 AOI22_X1 _08530_ (.A1(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[15][7] ),
    .A2(net111),
    .B1(net76),
    .B2(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[28][7] ),
    .ZN(_00209_));
 AOI22_X1 _08531_ (.A1(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[18][7] ),
    .A2(_00964_),
    .B1(net200),
    .B2(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[19][7] ),
    .ZN(_00210_));
 NAND4_X1 _08532_ (.A1(_00207_),
    .A2(_00208_),
    .A3(_00209_),
    .A4(_00210_),
    .ZN(_00211_));
 AOI22_X1 _08533_ (.A1(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[14][7] ),
    .A2(net88),
    .B1(net262),
    .B2(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[1][7] ),
    .ZN(_00212_));
 AOI22_X1 _08534_ (.A1(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[20][7] ),
    .A2(net246),
    .B1(_01007_),
    .B2(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[13][7] ),
    .ZN(_00213_));
 AOI22_X1 _08535_ (.A1(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[17][7] ),
    .A2(net81),
    .B1(_00996_),
    .B2(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[22][7] ),
    .ZN(_00214_));
 AOI22_X2 _08536_ (.A1(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[3][7] ),
    .A2(net63),
    .B1(_00993_),
    .B2(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[11][7] ),
    .ZN(_00215_));
 NAND4_X2 _08537_ (.A1(_00212_),
    .A2(_00213_),
    .A3(_00214_),
    .A4(_00215_),
    .ZN(_00216_));
 NOR4_X2 _08538_ (.A1(_00201_),
    .A2(_00206_),
    .A3(_00211_),
    .A4(_00216_),
    .ZN(_00217_));
 OAI21_X1 _08539_ (.A(_01662_),
    .B1(net130),
    .B2(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[0][7] ),
    .ZN(_00218_));
 OAI21_X1 _08540_ (.A(_01406_),
    .B1(_00217_),
    .B2(_00218_),
    .ZN(_00219_));
 NOR3_X1 _08541_ (.A1(_00151_),
    .A2(_00196_),
    .A3(_00219_),
    .ZN(_00220_));
 AOI22_X1 _08542_ (.A1(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[26][7] ),
    .A2(net169),
    .B1(net205),
    .B2(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[13][7] ),
    .ZN(_00221_));
 AOI22_X1 _08543_ (.A1(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[27][7] ),
    .A2(net189),
    .B1(net125),
    .B2(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[4][7] ),
    .ZN(_00222_));
 AND2_X1 _08544_ (.A1(_00221_),
    .A2(_00222_),
    .ZN(_00223_));
 AOI22_X1 _08545_ (.A1(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[24][7] ),
    .A2(net72),
    .B1(net85),
    .B2(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[14][7] ),
    .ZN(_00224_));
 AOI22_X1 _08546_ (.A1(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[17][7] ),
    .A2(net80),
    .B1(net67),
    .B2(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[7][7] ),
    .ZN(_00225_));
 AOI22_X1 _08547_ (.A1(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[18][7] ),
    .A2(net264),
    .B1(net247),
    .B2(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[20][7] ),
    .ZN(_00226_));
 AOI22_X1 _08548_ (.A1(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[8][7] ),
    .A2(net184),
    .B1(net210),
    .B2(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[30][7] ),
    .ZN(_00227_));
 AOI22_X1 _08549_ (.A1(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[1][7] ),
    .A2(net257),
    .B1(net197),
    .B2(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[19][7] ),
    .ZN(_00228_));
 AOI21_X1 _08550_ (.A(net113),
    .B1(net138),
    .B2(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[5][7] ),
    .ZN(_00229_));
 AND4_X1 _08551_ (.A1(_00226_),
    .A2(_00227_),
    .A3(_00228_),
    .A4(_00229_),
    .ZN(_00230_));
 AND4_X1 _08552_ (.A1(_00223_),
    .A2(_00224_),
    .A3(_00225_),
    .A4(_00230_),
    .ZN(_00231_));
 AOI22_X1 _08553_ (.A1(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[28][7] ),
    .A2(net75),
    .B1(net225),
    .B2(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[22][7] ),
    .ZN(_00232_));
 AOI22_X1 _08554_ (.A1(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[3][7] ),
    .A2(net64),
    .B1(net219),
    .B2(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[9][7] ),
    .ZN(_00233_));
 AND2_X1 _08555_ (.A1(_00232_),
    .A2(_00233_),
    .ZN(_00234_));
 AOI22_X1 _08556_ (.A1(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[6][7] ),
    .A2(net161),
    .B1(net154),
    .B2(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[25][7] ),
    .ZN(_00235_));
 AOI22_X1 _08557_ (.A1(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[29][7] ),
    .A2(net143),
    .B1(net234),
    .B2(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[11][7] ),
    .ZN(_00236_));
 AND2_X1 _08558_ (.A1(_00235_),
    .A2(_00236_),
    .ZN(_00237_));
 AOI22_X1 _08559_ (.A1(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[12][7] ),
    .A2(net270),
    .B1(net241),
    .B2(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[2][7] ),
    .ZN(_00238_));
 AOI22_X1 _08560_ (.A1(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[15][7] ),
    .A2(net106),
    .B1(net96),
    .B2(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[31][7] ),
    .ZN(_00239_));
 AOI22_X1 _08561_ (.A1(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[23][7] ),
    .A2(net105),
    .B1(net118),
    .B2(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[16][7] ),
    .ZN(_00240_));
 AOI22_X1 _08562_ (.A1(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[10][7] ),
    .A2(net91),
    .B1(net82),
    .B2(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[21][7] ),
    .ZN(_00241_));
 AND4_X1 _08563_ (.A1(_00238_),
    .A2(_00239_),
    .A3(_00240_),
    .A4(_00241_),
    .ZN(_00242_));
 AND4_X1 _08564_ (.A1(_00231_),
    .A2(_00234_),
    .A3(_00237_),
    .A4(_00242_),
    .ZN(_00243_));
 OAI21_X1 _08565_ (.A(_01350_),
    .B1(net130),
    .B2(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[0][7] ),
    .ZN(_00244_));
 AOI22_X1 _08566_ (.A1(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[23][7] ),
    .A2(net99),
    .B1(net253),
    .B2(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[1][7] ),
    .ZN(_00245_));
 AOI22_X1 _08567_ (.A1(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[12][7] ),
    .A2(net274),
    .B1(net206),
    .B2(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[13][7] ),
    .ZN(_00246_));
 AOI22_X1 _08568_ (.A1(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[16][7] ),
    .A2(net121),
    .B1(net150),
    .B2(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[25][7] ),
    .ZN(_00247_));
 AOI22_X1 _08569_ (.A1(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[29][7] ),
    .A2(net146),
    .B1(net244),
    .B2(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[20][7] ),
    .ZN(_00248_));
 NAND4_X2 _08570_ (.A1(_00245_),
    .A2(_00246_),
    .A3(_00247_),
    .A4(_00248_),
    .ZN(_00249_));
 AOI22_X1 _08571_ (.A1(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[6][7] ),
    .A2(net156),
    .B1(net215),
    .B2(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[30][7] ),
    .ZN(_00250_));
 AOI22_X1 _08572_ (.A1(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[10][7] ),
    .A2(net89),
    .B1(_00971_),
    .B2(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[14][7] ),
    .ZN(_00251_));
 AOI22_X1 _08573_ (.A1(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[4][7] ),
    .A2(net128),
    .B1(_00999_),
    .B2(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[9][7] ),
    .ZN(_00252_));
 AOI21_X1 _08574_ (.A(net115),
    .B1(net231),
    .B2(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[11][7] ),
    .ZN(_00253_));
 NAND4_X2 _08575_ (.A1(_00250_),
    .A2(_00251_),
    .A3(_00252_),
    .A4(_00253_),
    .ZN(_00254_));
 AOI22_X1 _08576_ (.A1(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[28][7] ),
    .A2(_01032_),
    .B1(net228),
    .B2(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[22][7] ),
    .ZN(_00255_));
 AOI22_X1 _08577_ (.A1(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[17][7] ),
    .A2(net81),
    .B1(_00981_),
    .B2(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[21][7] ),
    .ZN(_00256_));
 AOI22_X1 _08578_ (.A1(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[3][7] ),
    .A2(net63),
    .B1(_01149_),
    .B2(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[31][7] ),
    .ZN(_00257_));
 AOI22_X1 _08579_ (.A1(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[24][7] ),
    .A2(net73),
    .B1(net201),
    .B2(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[19][7] ),
    .ZN(_00258_));
 NAND4_X2 _08580_ (.A1(_00255_),
    .A2(_00256_),
    .A3(_00257_),
    .A4(_00258_),
    .ZN(_00259_));
 AOI22_X1 _08581_ (.A1(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[15][7] ),
    .A2(net112),
    .B1(net264),
    .B2(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[18][7] ),
    .ZN(_00260_));
 AOI22_X1 _08582_ (.A1(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[8][7] ),
    .A2(net176),
    .B1(net172),
    .B2(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[26][7] ),
    .ZN(_00261_));
 AOI22_X1 _08583_ (.A1(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[7][7] ),
    .A2(net70),
    .B1(_00989_),
    .B2(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[2][7] ),
    .ZN(_00262_));
 AOI22_X2 _08584_ (.A1(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[27][7] ),
    .A2(net186),
    .B1(net135),
    .B2(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[5][7] ),
    .ZN(_00263_));
 NAND4_X2 _08585_ (.A1(_00260_),
    .A2(_00261_),
    .A3(_00262_),
    .A4(_00263_),
    .ZN(_00264_));
 NOR4_X4 _08586_ (.A1(_00249_),
    .A2(_00254_),
    .A3(_00259_),
    .A4(_00264_),
    .ZN(_00265_));
 OAI21_X1 _08587_ (.A(_01731_),
    .B1(net130),
    .B2(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[0][7] ),
    .ZN(_00266_));
 AOI22_X1 _08588_ (.A1(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[3][7] ),
    .A2(net64),
    .B1(net163),
    .B2(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[6][7] ),
    .ZN(_00267_));
 AOI22_X1 _08589_ (.A1(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[16][7] ),
    .A2(net117),
    .B1(net194),
    .B2(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[19][7] ),
    .ZN(_00268_));
 AOI22_X1 _08590_ (.A1(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[22][7] ),
    .A2(net226),
    .B1(net204),
    .B2(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[13][7] ),
    .ZN(_00269_));
 AOI22_X1 _08591_ (.A1(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[28][7] ),
    .A2(net77),
    .B1(net153),
    .B2(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[25][7] ),
    .ZN(_00270_));
 NAND4_X1 _08592_ (.A1(_00267_),
    .A2(_00268_),
    .A3(_00269_),
    .A4(_00270_),
    .ZN(_00271_));
 AOI22_X1 _08593_ (.A1(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[8][7] ),
    .A2(net179),
    .B1(net219),
    .B2(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[9][7] ),
    .ZN(_00272_));
 AOI22_X1 _08594_ (.A1(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[18][7] ),
    .A2(net265),
    .B1(net256),
    .B2(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[1][7] ),
    .ZN(_00273_));
 AOI22_X1 _08595_ (.A1(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[26][7] ),
    .A2(net170),
    .B1(net85),
    .B2(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[14][7] ),
    .ZN(_00274_));
 AOI21_X1 _08596_ (.A(net113),
    .B1(net241),
    .B2(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[2][7] ),
    .ZN(_00275_));
 NAND4_X2 _08597_ (.A1(_00272_),
    .A2(_00273_),
    .A3(_00274_),
    .A4(_00275_),
    .ZN(_00276_));
 AOI22_X1 _08598_ (.A1(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[15][7] ),
    .A2(net106),
    .B1(net209),
    .B2(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[30][7] ),
    .ZN(_00277_));
 AOI22_X1 _08599_ (.A1(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[4][7] ),
    .A2(net124),
    .B1(net90),
    .B2(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[10][7] ),
    .ZN(_00278_));
 AOI22_X1 _08600_ (.A1(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[27][7] ),
    .A2(net190),
    .B1(net234),
    .B2(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[11][7] ),
    .ZN(_00279_));
 AOI22_X2 _08601_ (.A1(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[17][7] ),
    .A2(net80),
    .B1(net82),
    .B2(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[21][7] ),
    .ZN(_00280_));
 NAND4_X2 _08602_ (.A1(_00277_),
    .A2(_00278_),
    .A3(_00279_),
    .A4(_00280_),
    .ZN(_00281_));
 AOI22_X1 _08603_ (.A1(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[12][7] ),
    .A2(net269),
    .B1(net251),
    .B2(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[20][7] ),
    .ZN(_00282_));
 AOI22_X1 _08604_ (.A1(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[24][7] ),
    .A2(net74),
    .B1(net68),
    .B2(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[7][7] ),
    .ZN(_00283_));
 AOI22_X1 _08605_ (.A1(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[5][7] ),
    .A2(net132),
    .B1(net95),
    .B2(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[31][7] ),
    .ZN(_00284_));
 AOI22_X1 _08606_ (.A1(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[23][7] ),
    .A2(net101),
    .B1(net142),
    .B2(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[29][7] ),
    .ZN(_00285_));
 NAND4_X1 _08607_ (.A1(_00282_),
    .A2(_00283_),
    .A3(_00284_),
    .A4(_00285_),
    .ZN(_00286_));
 NOR4_X2 _08608_ (.A1(_00271_),
    .A2(_00276_),
    .A3(_00281_),
    .A4(_00286_),
    .ZN(_00287_));
 OAI21_X1 _08609_ (.A(_01539_),
    .B1(net130),
    .B2(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[0][7] ),
    .ZN(_00288_));
 OAI222_X2 _08610_ (.A1(_00243_),
    .A2(_00244_),
    .B1(_00265_),
    .B2(_00266_),
    .C1(_00287_),
    .C2(_00288_),
    .ZN(_00289_));
 AOI22_X1 _08611_ (.A1(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[28][7] ),
    .A2(net75),
    .B1(net87),
    .B2(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[14][7] ),
    .ZN(_00290_));
 AOI22_X1 _08612_ (.A1(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[4][7] ),
    .A2(net128),
    .B1(net272),
    .B2(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[12][7] ),
    .ZN(_00291_));
 AOI22_X1 _08613_ (.A1(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[8][7] ),
    .A2(net183),
    .B1(net139),
    .B2(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[5][7] ),
    .ZN(_00292_));
 AOI22_X1 _08614_ (.A1(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[2][7] ),
    .A2(net243),
    .B1(_00999_),
    .B2(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[9][7] ),
    .ZN(_00293_));
 NAND4_X1 _08615_ (.A1(_00290_),
    .A2(_00291_),
    .A3(_00292_),
    .A4(_00293_),
    .ZN(_00294_));
 AOI22_X1 _08616_ (.A1(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[30][7] ),
    .A2(net211),
    .B1(net206),
    .B2(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[13][7] ),
    .ZN(_00295_));
 AOI22_X1 _08617_ (.A1(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[27][7] ),
    .A2(net192),
    .B1(net237),
    .B2(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[11][7] ),
    .ZN(_00296_));
 AOI22_X1 _08618_ (.A1(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[17][7] ),
    .A2(net78),
    .B1(net252),
    .B2(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[20][7] ),
    .ZN(_00297_));
 AOI21_X1 _08619_ (.A(_01119_),
    .B1(net73),
    .B2(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[24][7] ),
    .ZN(_00298_));
 NAND4_X1 _08620_ (.A1(_00295_),
    .A2(_00296_),
    .A3(_00297_),
    .A4(_00298_),
    .ZN(_00299_));
 AOI22_X1 _08621_ (.A1(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[18][7] ),
    .A2(net264),
    .B1(net198),
    .B2(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[19][7] ),
    .ZN(_00300_));
 AOI22_X1 _08622_ (.A1(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[10][7] ),
    .A2(net89),
    .B1(net228),
    .B2(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[22][7] ),
    .ZN(_00301_));
 AOI22_X1 _08623_ (.A1(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[7][7] ),
    .A2(net70),
    .B1(net253),
    .B2(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[1][7] ),
    .ZN(_00302_));
 AOI22_X2 _08624_ (.A1(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[25][7] ),
    .A2(net150),
    .B1(net146),
    .B2(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[29][7] ),
    .ZN(_00303_));
 NAND4_X2 _08625_ (.A1(_00300_),
    .A2(_00301_),
    .A3(_00302_),
    .A4(_00303_),
    .ZN(_00304_));
 AOI22_X1 _08626_ (.A1(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[16][7] ),
    .A2(net119),
    .B1(net109),
    .B2(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[15][7] ),
    .ZN(_00305_));
 AOI22_X1 _08627_ (.A1(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[3][7] ),
    .A2(net65),
    .B1(net84),
    .B2(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[21][7] ),
    .ZN(_00306_));
 AOI22_X1 _08628_ (.A1(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[26][7] ),
    .A2(net171),
    .B1(_01149_),
    .B2(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[31][7] ),
    .ZN(_00307_));
 AOI22_X2 _08629_ (.A1(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[23][7] ),
    .A2(net99),
    .B1(net160),
    .B2(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[6][7] ),
    .ZN(_00308_));
 NAND4_X2 _08630_ (.A1(_00305_),
    .A2(_00306_),
    .A3(_00307_),
    .A4(_00308_),
    .ZN(_00309_));
 NOR4_X2 _08631_ (.A1(_00294_),
    .A2(_00299_),
    .A3(_00304_),
    .A4(_00309_),
    .ZN(_00310_));
 OAI21_X1 _08632_ (.A(_01408_),
    .B1(net130),
    .B2(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[0][7] ),
    .ZN(_00311_));
 AOI22_X1 _08633_ (.A1(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[6][7] ),
    .A2(net158),
    .B1(net87),
    .B2(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[14][7] ),
    .ZN(_00312_));
 AOI22_X1 _08634_ (.A1(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[26][7] ),
    .A2(net174),
    .B1(net144),
    .B2(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[29][7] ),
    .ZN(_00313_));
 AOI22_X1 _08635_ (.A1(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[24][7] ),
    .A2(net71),
    .B1(net69),
    .B2(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[7][7] ),
    .ZN(_00314_));
 AOI22_X1 _08636_ (.A1(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[31][7] ),
    .A2(net93),
    .B1(net268),
    .B2(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[12][7] ),
    .ZN(_00315_));
 NAND4_X1 _08637_ (.A1(_00312_),
    .A2(_00313_),
    .A3(_00314_),
    .A4(_00315_),
    .ZN(_00316_));
 AOI22_X1 _08638_ (.A1(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[28][7] ),
    .A2(net76),
    .B1(net240),
    .B2(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[2][7] ),
    .ZN(_00317_));
 AOI22_X1 _08639_ (.A1(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[1][7] ),
    .A2(net254),
    .B1(net213),
    .B2(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[30][7] ),
    .ZN(_00318_));
 AOI22_X1 _08640_ (.A1(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[20][7] ),
    .A2(net245),
    .B1(net222),
    .B2(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[22][7] ),
    .ZN(_00319_));
 AOI21_X1 _08641_ (.A(net114),
    .B1(net196),
    .B2(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[19][7] ),
    .ZN(_00320_));
 NAND4_X2 _08642_ (.A1(_00317_),
    .A2(_00318_),
    .A3(_00319_),
    .A4(_00320_),
    .ZN(_00321_));
 AOI22_X1 _08643_ (.A1(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[21][7] ),
    .A2(net83),
    .B1(net229),
    .B2(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[11][7] ),
    .ZN(_00322_));
 AOI22_X1 _08644_ (.A1(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[8][7] ),
    .A2(net178),
    .B1(net217),
    .B2(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[9][7] ),
    .ZN(_00323_));
 AOI22_X1 _08645_ (.A1(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[17][7] ),
    .A2(net79),
    .B1(net188),
    .B2(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[27][7] ),
    .ZN(_00324_));
 AOI22_X2 _08646_ (.A1(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[18][7] ),
    .A2(net263),
    .B1(net203),
    .B2(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[13][7] ),
    .ZN(_00325_));
 NAND4_X2 _08647_ (.A1(_00322_),
    .A2(_00323_),
    .A3(_00324_),
    .A4(_00325_),
    .ZN(_00326_));
 AOI22_X1 _08648_ (.A1(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[16][7] ),
    .A2(net120),
    .B1(net126),
    .B2(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[4][7] ),
    .ZN(_00327_));
 AOI22_X1 _08649_ (.A1(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[3][7] ),
    .A2(net66),
    .B1(_00956_),
    .B2(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[10][7] ),
    .ZN(_00328_));
 AOI22_X1 _08650_ (.A1(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[23][7] ),
    .A2(net102),
    .B1(net134),
    .B2(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[5][7] ),
    .ZN(_00329_));
 AOI22_X1 _08651_ (.A1(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[15][7] ),
    .A2(net108),
    .B1(net148),
    .B2(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[25][7] ),
    .ZN(_00330_));
 NAND4_X1 _08652_ (.A1(_00327_),
    .A2(_00328_),
    .A3(_00329_),
    .A4(_00330_),
    .ZN(_00331_));
 NOR4_X2 _08653_ (.A1(_00316_),
    .A2(_00321_),
    .A3(_00326_),
    .A4(_00331_),
    .ZN(_00332_));
 OAI21_X1 _08654_ (.A(_01295_),
    .B1(net130),
    .B2(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[0][7] ),
    .ZN(_00333_));
 OAI22_X2 _08655_ (.A1(_00310_),
    .A2(_00311_),
    .B1(_00332_),
    .B2(_00333_),
    .ZN(_00334_));
 AOI22_X1 _08656_ (.A1(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[23][7] ),
    .A2(net98),
    .B1(net72),
    .B2(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[24][7] ),
    .ZN(_00335_));
 AOI22_X1 _08657_ (.A1(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[27][7] ),
    .A2(net191),
    .B1(net109),
    .B2(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[15][7] ),
    .ZN(_00336_));
 AOI22_X1 _08658_ (.A1(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[12][7] ),
    .A2(net266),
    .B1(net86),
    .B2(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[14][7] ),
    .ZN(_00337_));
 AOI22_X1 _08659_ (.A1(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[28][7] ),
    .A2(net75),
    .B1(net258),
    .B2(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[1][7] ),
    .ZN(_00338_));
 NAND4_X1 _08660_ (.A1(_00335_),
    .A2(_00336_),
    .A3(_00337_),
    .A4(_00338_),
    .ZN(_00339_));
 AOI22_X1 _08661_ (.A1(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[29][7] ),
    .A2(net145),
    .B1(net91),
    .B2(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[10][7] ),
    .ZN(_00340_));
 AOI22_X1 _08662_ (.A1(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[26][7] ),
    .A2(net168),
    .B1(net206),
    .B2(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[13][7] ),
    .ZN(_00341_));
 AOI22_X1 _08663_ (.A1(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[17][7] ),
    .A2(net78),
    .B1(net67),
    .B2(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[7][7] ),
    .ZN(_00342_));
 AOI21_X1 _08664_ (.A(net113),
    .B1(net164),
    .B2(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[6][7] ),
    .ZN(_00343_));
 NAND4_X1 _08665_ (.A1(_00340_),
    .A2(_00341_),
    .A3(_00342_),
    .A4(_00343_),
    .ZN(_00344_));
 AOI22_X1 _08666_ (.A1(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[3][7] ),
    .A2(net65),
    .B1(net128),
    .B2(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[4][7] ),
    .ZN(_00345_));
 AOI22_X1 _08667_ (.A1(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[16][7] ),
    .A2(net119),
    .B1(net220),
    .B2(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[9][7] ),
    .ZN(_00346_));
 AOI22_X1 _08668_ (.A1(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[5][7] ),
    .A2(net136),
    .B1(net207),
    .B2(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[30][7] ),
    .ZN(_00347_));
 AOI22_X1 _08669_ (.A1(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[21][7] ),
    .A2(net84),
    .B1(net232),
    .B2(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[11][7] ),
    .ZN(_00348_));
 NAND4_X1 _08670_ (.A1(_00345_),
    .A2(_00346_),
    .A3(_00347_),
    .A4(_00348_),
    .ZN(_00349_));
 AOI22_X1 _08671_ (.A1(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[8][7] ),
    .A2(net182),
    .B1(net198),
    .B2(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[19][7] ),
    .ZN(_00350_));
 AOI22_X1 _08672_ (.A1(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[18][7] ),
    .A2(net264),
    .B1(net248),
    .B2(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[20][7] ),
    .ZN(_00351_));
 AOI22_X1 _08673_ (.A1(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[25][7] ),
    .A2(net149),
    .B1(net243),
    .B2(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[2][7] ),
    .ZN(_00352_));
 AOI22_X2 _08674_ (.A1(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[31][7] ),
    .A2(_01149_),
    .B1(net223),
    .B2(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[22][7] ),
    .ZN(_00353_));
 NAND4_X2 _08675_ (.A1(_00350_),
    .A2(_00351_),
    .A3(_00352_),
    .A4(_00353_),
    .ZN(_00354_));
 NOR4_X2 _08676_ (.A1(_00339_),
    .A2(_00344_),
    .A3(_00349_),
    .A4(_00354_),
    .ZN(_00355_));
 OAI21_X1 _08677_ (.A(_00923_),
    .B1(net130),
    .B2(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[0][7] ),
    .ZN(_00356_));
 AOI22_X1 _08678_ (.A1(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[17][7] ),
    .A2(net80),
    .B1(net64),
    .B2(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[3][7] ),
    .ZN(_00357_));
 AOI22_X1 _08679_ (.A1(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[21][7] ),
    .A2(net83),
    .B1(net251),
    .B2(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[20][7] ),
    .ZN(_00358_));
 AOI22_X1 _08680_ (.A1(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[12][7] ),
    .A2(net269),
    .B1(net87),
    .B2(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[14][7] ),
    .ZN(_00359_));
 AOI22_X1 _08681_ (.A1(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[27][7] ),
    .A2(net192),
    .B1(net212),
    .B2(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[30][7] ),
    .ZN(_00360_));
 NAND4_X1 _08682_ (.A1(_00357_),
    .A2(_00358_),
    .A3(_00359_),
    .A4(_00360_),
    .ZN(_00361_));
 AOI22_X1 _08683_ (.A1(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[28][7] ),
    .A2(net77),
    .B1(net181),
    .B2(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[8][7] ),
    .ZN(_00362_));
 AOI22_X1 _08684_ (.A1(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[29][7] ),
    .A2(net144),
    .B1(net71),
    .B2(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[24][7] ),
    .ZN(_00363_));
 AOI22_X1 _08685_ (.A1(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[7][7] ),
    .A2(net68),
    .B1(net93),
    .B2(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[31][7] ),
    .ZN(_00364_));
 AOI21_X1 _08686_ (.A(net114),
    .B1(net263),
    .B2(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[18][7] ),
    .ZN(_00365_));
 NAND4_X1 _08687_ (.A1(_00362_),
    .A2(_00363_),
    .A3(_00364_),
    .A4(_00365_),
    .ZN(_00366_));
 AOI22_X1 _08688_ (.A1(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[6][7] ),
    .A2(net163),
    .B1(net193),
    .B2(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[19][7] ),
    .ZN(_00367_));
 AOI22_X1 _08689_ (.A1(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[23][7] ),
    .A2(net104),
    .B1(net260),
    .B2(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[1][7] ),
    .ZN(_00368_));
 AOI22_X1 _08690_ (.A1(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[16][7] ),
    .A2(net116),
    .B1(net132),
    .B2(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[5][7] ),
    .ZN(_00369_));
 AOI22_X1 _08691_ (.A1(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[15][7] ),
    .A2(net108),
    .B1(net217),
    .B2(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[9][7] ),
    .ZN(_00370_));
 NAND4_X1 _08692_ (.A1(_00367_),
    .A2(_00368_),
    .A3(_00369_),
    .A4(_00370_),
    .ZN(_00371_));
 AOI22_X1 _08693_ (.A1(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[2][7] ),
    .A2(net240),
    .B1(net236),
    .B2(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[11][7] ),
    .ZN(_00372_));
 AOI22_X1 _08694_ (.A1(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[26][7] ),
    .A2(net175),
    .B1(net222),
    .B2(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[22][7] ),
    .ZN(_00373_));
 AOI22_X1 _08695_ (.A1(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[25][7] ),
    .A2(net148),
    .B1(net126),
    .B2(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[4][7] ),
    .ZN(_00374_));
 AOI22_X1 _08696_ (.A1(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[10][7] ),
    .A2(net90),
    .B1(net203),
    .B2(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[13][7] ),
    .ZN(_00375_));
 NAND4_X1 _08697_ (.A1(_00372_),
    .A2(_00373_),
    .A3(_00374_),
    .A4(_00375_),
    .ZN(_00376_));
 NOR4_X1 _08698_ (.A1(_00361_),
    .A2(_00366_),
    .A3(_00371_),
    .A4(_00376_),
    .ZN(_00377_));
 OAI21_X1 _08699_ (.A(_01700_),
    .B1(net130),
    .B2(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[0][7] ),
    .ZN(_00378_));
 OAI22_X1 _08700_ (.A1(_00355_),
    .A2(_00356_),
    .B1(_00377_),
    .B2(_00378_),
    .ZN(_00379_));
 INV_X1 _08701_ (.A(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[8][7] ),
    .ZN(_00380_));
 OAI21_X1 _08702_ (.A(net130),
    .B1(_03001_),
    .B2(_00380_),
    .ZN(_00381_));
 AOI221_X2 _08703_ (.A(_00381_),
    .B1(net157),
    .B2(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[6][7] ),
    .C1(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[23][7] ),
    .C2(net102),
    .ZN(_00382_));
 INV_X1 _08704_ (.A(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[16][7] ),
    .ZN(_00383_));
 INV_X1 _08705_ (.A(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[20][7] ),
    .ZN(_00384_));
 OAI22_X1 _08706_ (.A1(_00383_),
    .A2(_01027_),
    .B1(_01691_),
    .B2(_00384_),
    .ZN(_00385_));
 AOI221_X2 _08707_ (.A(_00385_),
    .B1(_01102_),
    .B2(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[3][7] ),
    .C1(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[24][7] ),
    .C2(_01059_),
    .ZN(_00386_));
 INV_X1 _08708_ (.A(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[29][7] ),
    .ZN(_00387_));
 INV_X1 _08709_ (.A(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[2][7] ),
    .ZN(_00388_));
 OAI22_X1 _08710_ (.A1(_00387_),
    .A2(_01425_),
    .B1(_01211_),
    .B2(_00388_),
    .ZN(_00389_));
 AOI221_X2 _08711_ (.A(_00389_),
    .B1(net69),
    .B2(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[7][7] ),
    .C1(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[12][7] ),
    .C2(_00950_),
    .ZN(_00390_));
 AOI22_X1 _08712_ (.A1(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[27][7] ),
    .A2(net187),
    .B1(net199),
    .B2(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[19][7] ),
    .ZN(_00391_));
 AOI22_X1 _08713_ (.A1(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[5][7] ),
    .A2(net133),
    .B1(net203),
    .B2(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[13][7] ),
    .ZN(_00392_));
 AND2_X1 _08714_ (.A1(_00391_),
    .A2(_00392_),
    .ZN(_00393_));
 NAND4_X2 _08715_ (.A1(_00382_),
    .A2(_00386_),
    .A3(_00390_),
    .A4(_00393_),
    .ZN(_00394_));
 INV_X1 _08716_ (.A(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[15][7] ),
    .ZN(_00395_));
 INV_X1 _08717_ (.A(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[22][7] ),
    .ZN(_00396_));
 OAI22_X1 _08718_ (.A1(_00395_),
    .A2(_01029_),
    .B1(_01216_),
    .B2(_00396_),
    .ZN(_00397_));
 AOI221_X2 _08719_ (.A(_00397_),
    .B1(net174),
    .B2(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[26][7] ),
    .C1(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[28][7] ),
    .C2(net76),
    .ZN(_00398_));
 INV_X1 _08720_ (.A(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[25][7] ),
    .ZN(_00399_));
 INV_X1 _08721_ (.A(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[4][7] ),
    .ZN(_00400_));
 OAI22_X2 _08722_ (.A1(_00399_),
    .A2(_01470_),
    .B1(_00941_),
    .B2(_00400_),
    .ZN(_00401_));
 AOI221_X2 _08723_ (.A(_00401_),
    .B1(net229),
    .B2(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[11][7] ),
    .C1(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[21][7] ),
    .C2(net83),
    .ZN(_00402_));
 INV_X1 _08724_ (.A(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[18][7] ),
    .ZN(_00403_));
 INV_X1 _08725_ (.A(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[1][7] ),
    .ZN(_00404_));
 OAI22_X2 _08726_ (.A1(_00403_),
    .A2(_02024_),
    .B1(_01210_),
    .B2(_00404_),
    .ZN(_00405_));
 AOI221_X2 _08727_ (.A(_00405_),
    .B1(net88),
    .B2(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[14][7] ),
    .C1(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[17][7] ),
    .C2(net81),
    .ZN(_00406_));
 INV_X1 _08728_ (.A(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[31][7] ),
    .ZN(_00407_));
 INV_X1 _08729_ (.A(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[9][7] ),
    .ZN(_00408_));
 OAI22_X1 _08730_ (.A1(_00407_),
    .A2(_00934_),
    .B1(_01420_),
    .B2(_00408_),
    .ZN(_00409_));
 AOI221_X2 _08731_ (.A(_00409_),
    .B1(_00956_),
    .B2(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[10][7] ),
    .C1(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[30][7] ),
    .C2(net213),
    .ZN(_00410_));
 NAND4_X2 _08732_ (.A1(_00398_),
    .A2(_00402_),
    .A3(_00406_),
    .A4(_00410_),
    .ZN(_00411_));
 OAI221_X2 _08733_ (.A(_01583_),
    .B1(_00394_),
    .B2(_00411_),
    .C1(net130),
    .C2(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[0][7] ),
    .ZN(_00412_));
 AOI22_X1 _08734_ (.A1(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[16][7] ),
    .A2(net121),
    .B1(net274),
    .B2(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[12][7] ),
    .ZN(_00413_));
 AOI22_X1 _08735_ (.A1(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[1][7] ),
    .A2(net262),
    .B1(net215),
    .B2(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[30][7] ),
    .ZN(_00414_));
 AND2_X1 _08736_ (.A1(_00413_),
    .A2(_00414_),
    .ZN(_00415_));
 INV_X1 _08737_ (.A(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[28][7] ),
    .ZN(_00416_));
 NAND2_X1 _08738_ (.A1(net9),
    .A2(_00937_),
    .ZN(_00417_));
 INV_X1 _08739_ (.A(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[6][7] ),
    .ZN(_00418_));
 OAI33_X1 _08740_ (.A1(_00416_),
    .A2(_00979_),
    .A3(_00970_),
    .B1(_00417_),
    .B2(_00952_),
    .B3(_00418_),
    .ZN(_00419_));
 AOI221_X2 _08741_ (.A(_00419_),
    .B1(net88),
    .B2(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[14][7] ),
    .C1(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[21][7] ),
    .C2(_00981_),
    .ZN(_00420_));
 INV_X1 _08742_ (.A(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[15][7] ),
    .ZN(_00421_));
 INV_X1 _08743_ (.A(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[13][7] ),
    .ZN(_00422_));
 OAI22_X2 _08744_ (.A1(_00421_),
    .A2(_01029_),
    .B1(_03431_),
    .B2(_00422_),
    .ZN(_00423_));
 AOI221_X2 _08745_ (.A(_00423_),
    .B1(net63),
    .B2(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[3][7] ),
    .C1(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[29][7] ),
    .C2(_01050_),
    .ZN(_00424_));
 INV_X1 _08746_ (.A(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[31][7] ),
    .ZN(_00425_));
 INV_X1 _08747_ (.A(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[2][7] ),
    .ZN(_00426_));
 OAI22_X1 _08748_ (.A1(_00425_),
    .A2(_00934_),
    .B1(_01211_),
    .B2(_00426_),
    .ZN(_00427_));
 AOI221_X2 _08749_ (.A(_00427_),
    .B1(net89),
    .B2(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[10][7] ),
    .C1(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[26][7] ),
    .C2(net172),
    .ZN(_00428_));
 NAND4_X2 _08750_ (.A1(_00415_),
    .A2(_00420_),
    .A3(_00424_),
    .A4(_00428_),
    .ZN(_00429_));
 NAND3_X1 _08751_ (.A1(net8),
    .A2(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[11][7] ),
    .A3(_01418_),
    .ZN(_00430_));
 OAI21_X1 _08752_ (.A(_00430_),
    .B1(_00985_),
    .B2(net8),
    .ZN(_00431_));
 AOI222_X2 _08753_ (.A1(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[17][7] ),
    .A2(net81),
    .B1(_03867_),
    .B2(_00431_),
    .C1(net129),
    .C2(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[4][7] ),
    .ZN(_00432_));
 INV_X1 _08754_ (.A(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[8][7] ),
    .ZN(_00433_));
 INV_X1 _08755_ (.A(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[18][7] ),
    .ZN(_00434_));
 OAI22_X1 _08756_ (.A1(_00433_),
    .A2(_03001_),
    .B1(_02024_),
    .B2(_00434_),
    .ZN(_00435_));
 AOI221_X2 _08757_ (.A(_00435_),
    .B1(net73),
    .B2(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[24][7] ),
    .C1(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[27][7] ),
    .C2(net186),
    .ZN(_00436_));
 AOI22_X1 _08758_ (.A1(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[5][7] ),
    .A2(_01057_),
    .B1(_00986_),
    .B2(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[20][7] ),
    .ZN(_00437_));
 AOI22_X1 _08759_ (.A1(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[9][7] ),
    .A2(net221),
    .B1(net201),
    .B2(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[19][7] ),
    .ZN(_00438_));
 AND2_X1 _08760_ (.A1(_00437_),
    .A2(_00438_),
    .ZN(_00439_));
 INV_X1 _08761_ (.A(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[23][7] ),
    .ZN(_00440_));
 INV_X1 _08762_ (.A(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[25][7] ),
    .ZN(_00441_));
 OAI22_X1 _08763_ (.A1(_00440_),
    .A2(_01417_),
    .B1(_01470_),
    .B2(_00441_),
    .ZN(_00442_));
 AOI221_X2 _08764_ (.A(_00442_),
    .B1(net70),
    .B2(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[7][7] ),
    .C1(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[22][7] ),
    .C2(net228),
    .ZN(_00443_));
 NAND4_X2 _08765_ (.A1(_00432_),
    .A2(_00436_),
    .A3(_00439_),
    .A4(_00443_),
    .ZN(_00444_));
 OAI221_X2 _08766_ (.A(_01502_),
    .B1(_00429_),
    .B2(_00444_),
    .C1(_01064_),
    .C2(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[0][7] ),
    .ZN(_00445_));
 AND3_X1 _08767_ (.A1(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[3][7] ),
    .A2(_02035_),
    .A3(_02036_),
    .ZN(_00446_));
 AND3_X1 _08768_ (.A1(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[24][7] ),
    .A2(_01121_),
    .A3(_02912_),
    .ZN(_00447_));
 INV_X1 _08769_ (.A(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[15][7] ),
    .ZN(_00448_));
 INV_X1 _08770_ (.A(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[26][7] ),
    .ZN(_00449_));
 OAI22_X1 _08771_ (.A1(_00448_),
    .A2(_01029_),
    .B1(_01203_),
    .B2(_00449_),
    .ZN(_00450_));
 NOR4_X1 _08772_ (.A1(net114),
    .A2(_00446_),
    .A3(_00447_),
    .A4(_00450_),
    .ZN(_00451_));
 INV_X1 _08773_ (.A(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[2][7] ),
    .ZN(_00452_));
 INV_X1 _08774_ (.A(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[22][7] ),
    .ZN(_00453_));
 OAI22_X1 _08775_ (.A1(_00452_),
    .A2(_01211_),
    .B1(_01216_),
    .B2(_00453_),
    .ZN(_00454_));
 AOI221_X1 _08776_ (.A(_00454_),
    .B1(net138),
    .B2(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[5][7] ),
    .C1(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[21][7] ),
    .C2(net83),
    .ZN(_00455_));
 INV_X1 _08777_ (.A(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[20][7] ),
    .ZN(_00456_));
 INV_X1 _08778_ (.A(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[19][7] ),
    .ZN(_00457_));
 OAI22_X1 _08779_ (.A1(_00456_),
    .A2(_01691_),
    .B1(_03436_),
    .B2(_00457_),
    .ZN(_00458_));
 AOI221_X1 _08780_ (.A(_00458_),
    .B1(net126),
    .B2(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[4][7] ),
    .C1(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[28][7] ),
    .C2(net77),
    .ZN(_00459_));
 INV_X1 _08781_ (.A(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[9][7] ),
    .ZN(_00460_));
 INV_X1 _08782_ (.A(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[30][7] ),
    .ZN(_00461_));
 OAI22_X1 _08783_ (.A1(_00460_),
    .A2(_01420_),
    .B1(_01204_),
    .B2(_00461_),
    .ZN(_00462_));
 AOI221_X2 _08784_ (.A(_00462_),
    .B1(net86),
    .B2(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[14][7] ),
    .C1(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[29][7] ),
    .C2(net143),
    .ZN(_00463_));
 NAND4_X1 _08785_ (.A1(_00451_),
    .A2(_00455_),
    .A3(_00459_),
    .A4(_00463_),
    .ZN(_00464_));
 AOI22_X1 _08786_ (.A1(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[23][7] ),
    .A2(net104),
    .B1(net164),
    .B2(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[6][7] ),
    .ZN(_00465_));
 AOI22_X1 _08787_ (.A1(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[17][7] ),
    .A2(net78),
    .B1(_01076_),
    .B2(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[7][7] ),
    .ZN(_00466_));
 INV_X1 _08788_ (.A(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[1][7] ),
    .ZN(_00467_));
 INV_X1 _08789_ (.A(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[11][7] ),
    .ZN(_00468_));
 OAI22_X1 _08790_ (.A1(_00467_),
    .A2(_01210_),
    .B1(_02556_),
    .B2(_00468_),
    .ZN(_00469_));
 AOI221_X1 _08791_ (.A(_00469_),
    .B1(net91),
    .B2(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[10][7] ),
    .C1(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[16][7] ),
    .C2(_01097_),
    .ZN(_00470_));
 AOI22_X1 _08792_ (.A1(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[27][7] ),
    .A2(net192),
    .B1(net181),
    .B2(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[8][7] ),
    .ZN(_00471_));
 AOI222_X2 _08793_ (.A1(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[25][7] ),
    .A2(_01046_),
    .B1(net205),
    .B2(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[13][7] ),
    .C1(net95),
    .C2(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[31][7] ),
    .ZN(_00472_));
 AOI22_X1 _08794_ (.A1(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[12][7] ),
    .A2(_00950_),
    .B1(net263),
    .B2(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[18][7] ),
    .ZN(_00473_));
 AND3_X1 _08795_ (.A1(_00471_),
    .A2(_00472_),
    .A3(_00473_),
    .ZN(_00474_));
 NAND4_X1 _08796_ (.A1(_00465_),
    .A2(_00466_),
    .A3(_00470_),
    .A4(_00474_),
    .ZN(_00475_));
 OAI221_X2 _08797_ (.A(_01764_),
    .B1(_00464_),
    .B2(_00475_),
    .C1(net130),
    .C2(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[0][7] ),
    .ZN(_00476_));
 INV_X1 _08798_ (.A(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[27][7] ),
    .ZN(_00477_));
 INV_X1 _08799_ (.A(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[31][7] ),
    .ZN(_00478_));
 OAI22_X1 _08800_ (.A1(_00477_),
    .A2(_02555_),
    .B1(_00934_),
    .B2(_00478_),
    .ZN(_00479_));
 AOI221_X1 _08801_ (.A(_00479_),
    .B1(_01102_),
    .B2(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[3][7] ),
    .C1(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[11][7] ),
    .C2(net229),
    .ZN(_00480_));
 MUX2_X1 _08802_ (.A(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[12][7] ),
    .B(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[14][7] ),
    .S(net8),
    .Z(_00481_));
 AOI221_X2 _08803_ (.A(net115),
    .B1(net92),
    .B2(_00481_),
    .C1(net148),
    .C2(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[25][7] ),
    .ZN(_00482_));
 AOI22_X1 _08804_ (.A1(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[1][7] ),
    .A2(net261),
    .B1(net227),
    .B2(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[22][7] ),
    .ZN(_00483_));
 AOI22_X1 _08805_ (.A1(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[13][7] ),
    .A2(net203),
    .B1(net202),
    .B2(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[19][7] ),
    .ZN(_00484_));
 AND2_X1 _08806_ (.A1(_00483_),
    .A2(_00484_),
    .ZN(_00485_));
 INV_X1 _08807_ (.A(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[17][7] ),
    .ZN(_00486_));
 INV_X1 _08808_ (.A(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[23][7] ),
    .ZN(_00487_));
 OAI33_X1 _08809_ (.A1(_00486_),
    .A2(_01015_),
    .A3(_00979_),
    .B1(_00960_),
    .B2(_00980_),
    .B3(_00487_),
    .ZN(_00488_));
 AOI221_X2 _08810_ (.A(_00488_),
    .B1(net158),
    .B2(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[6][7] ),
    .C1(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[10][7] ),
    .C2(_00956_),
    .ZN(_00489_));
 NAND4_X2 _08811_ (.A1(_00480_),
    .A2(_00482_),
    .A3(_00485_),
    .A4(_00489_),
    .ZN(_00490_));
 INV_X1 _08812_ (.A(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[18][7] ),
    .ZN(_00491_));
 INV_X1 _08813_ (.A(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[2][7] ),
    .ZN(_00492_));
 OAI22_X1 _08814_ (.A1(_00491_),
    .A2(_02024_),
    .B1(_01211_),
    .B2(_00492_),
    .ZN(_00493_));
 AOI221_X1 _08815_ (.A(_00493_),
    .B1(net69),
    .B2(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[7][7] ),
    .C1(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[16][7] ),
    .C2(net122),
    .ZN(_00494_));
 INV_X1 _08816_ (.A(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[5][7] ),
    .ZN(_00495_));
 INV_X1 _08817_ (.A(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[9][7] ),
    .ZN(_00496_));
 OAI22_X1 _08818_ (.A1(_00495_),
    .A2(_02238_),
    .B1(_01420_),
    .B2(_00496_),
    .ZN(_00497_));
 AOI221_X1 _08819_ (.A(_00497_),
    .B1(net245),
    .B2(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[20][7] ),
    .C1(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[28][7] ),
    .C2(net76),
    .ZN(_00498_));
 AOI22_X1 _08820_ (.A1(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[26][7] ),
    .A2(_01038_),
    .B1(net126),
    .B2(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[4][7] ),
    .ZN(_00499_));
 AOI22_X1 _08821_ (.A1(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[15][7] ),
    .A2(net111),
    .B1(net214),
    .B2(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[30][7] ),
    .ZN(_00500_));
 AND2_X1 _08822_ (.A1(_00499_),
    .A2(_00500_),
    .ZN(_00501_));
 INV_X1 _08823_ (.A(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[21][7] ),
    .ZN(_00502_));
 INV_X1 _08824_ (.A(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[8][7] ),
    .ZN(_00503_));
 OAI33_X1 _08825_ (.A1(_00502_),
    .A2(_00979_),
    .A3(_00980_),
    .B1(_00948_),
    .B2(_00954_),
    .B3(_00503_),
    .ZN(_00504_));
 AOI221_X1 _08826_ (.A(_00504_),
    .B1(_01059_),
    .B2(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[24][7] ),
    .C1(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[29][7] ),
    .C2(net141),
    .ZN(_00505_));
 NAND4_X1 _08827_ (.A1(_00494_),
    .A2(_00498_),
    .A3(_00501_),
    .A4(_00505_),
    .ZN(_00506_));
 OAI221_X2 _08828_ (.A(_01623_),
    .B1(_00490_),
    .B2(_00506_),
    .C1(net130),
    .C2(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[0][7] ),
    .ZN(_00507_));
 NAND4_X2 _08829_ (.A1(_00412_),
    .A2(_00445_),
    .A3(_00476_),
    .A4(_00507_),
    .ZN(_00508_));
 NOR4_X2 _08830_ (.A1(_00289_),
    .A2(_00334_),
    .A3(_00379_),
    .A4(_00508_),
    .ZN(_00509_));
 AOI22_X1 _08831_ (.A1(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[1][7] ),
    .A2(net256),
    .B1(net217),
    .B2(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[9][7] ),
    .ZN(_00510_));
 AOI22_X1 _08832_ (.A1(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[14][7] ),
    .A2(net85),
    .B1(net82),
    .B2(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[21][7] ),
    .ZN(_00511_));
 AOI22_X1 _08833_ (.A1(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[17][7] ),
    .A2(net79),
    .B1(net132),
    .B2(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[5][7] ),
    .ZN(_00512_));
 AOI22_X1 _08834_ (.A1(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[28][7] ),
    .A2(net77),
    .B1(net173),
    .B2(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[26][7] ),
    .ZN(_00513_));
 NAND4_X1 _08835_ (.A1(_00510_),
    .A2(_00511_),
    .A3(_00512_),
    .A4(_00513_),
    .ZN(_00514_));
 AOI22_X1 _08836_ (.A1(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[23][7] ),
    .A2(net100),
    .B1(net95),
    .B2(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[31][7] ),
    .ZN(_00515_));
 AOI22_X1 _08837_ (.A1(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[25][7] ),
    .A2(net153),
    .B1(net74),
    .B2(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[24][7] ),
    .ZN(_00516_));
 AOI22_X1 _08838_ (.A1(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[15][7] ),
    .A2(net107),
    .B1(net204),
    .B2(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[13][7] ),
    .ZN(_00517_));
 AOI21_X1 _08839_ (.A(net113),
    .B1(net64),
    .B2(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[3][7] ),
    .ZN(_00518_));
 NAND4_X1 _08840_ (.A1(_00515_),
    .A2(_00516_),
    .A3(_00517_),
    .A4(_00518_),
    .ZN(_00519_));
 AOI22_X1 _08841_ (.A1(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[8][7] ),
    .A2(net181),
    .B1(net263),
    .B2(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[18][7] ),
    .ZN(_00520_));
 AOI22_X1 _08842_ (.A1(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[6][7] ),
    .A2(net162),
    .B1(net208),
    .B2(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[30][7] ),
    .ZN(_00521_));
 AOI22_X1 _08843_ (.A1(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[29][7] ),
    .A2(net142),
    .B1(net267),
    .B2(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[12][7] ),
    .ZN(_00522_));
 AOI22_X1 _08844_ (.A1(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[7][7] ),
    .A2(net68),
    .B1(net250),
    .B2(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[20][7] ),
    .ZN(_00523_));
 NAND4_X1 _08845_ (.A1(_00520_),
    .A2(_00521_),
    .A3(_00522_),
    .A4(_00523_),
    .ZN(_00524_));
 AOI22_X1 _08846_ (.A1(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[10][7] ),
    .A2(net90),
    .B1(net242),
    .B2(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[2][7] ),
    .ZN(_00525_));
 AOI22_X1 _08847_ (.A1(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[16][7] ),
    .A2(net116),
    .B1(net226),
    .B2(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[22][7] ),
    .ZN(_00526_));
 AOI22_X1 _08848_ (.A1(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[27][7] ),
    .A2(net190),
    .B1(net194),
    .B2(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[19][7] ),
    .ZN(_00527_));
 AOI22_X1 _08849_ (.A1(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[4][7] ),
    .A2(net123),
    .B1(net233),
    .B2(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[11][7] ),
    .ZN(_00528_));
 NAND4_X1 _08850_ (.A1(_00525_),
    .A2(_00526_),
    .A3(_00527_),
    .A4(_00528_),
    .ZN(_00529_));
 OR4_X2 _08851_ (.A1(_00514_),
    .A2(_00519_),
    .A3(_00524_),
    .A4(_00529_),
    .ZN(_00530_));
 OAI21_X1 _08852_ (.A(_00530_),
    .B1(net130),
    .B2(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[0][7] ),
    .ZN(_00531_));
 AOI221_X2 _08853_ (.A(_00907_),
    .B1(_00220_),
    .B2(_00509_),
    .C1(_00531_),
    .C2(_01820_),
    .ZN(\rdata_o_n[7] ));
 AND2_X1 _08854_ (.A1(\lut.cg_we_global.clk_en ),
    .A2(clknet_3_0__leaf_clk_i),
    .ZN(_00532_));
 TAPCELL_X1 PHY_56 ();
 TAPCELL_X1 PHY_55 ();
 AND2_X1 _08857_ (.A1(\lut.gen_sub_units_scm.__15.sub_unit_i.cg_we_global.clk_en ),
    .A2(clknet_2_2__leaf__00532_),
    .ZN(_00534_));
 TAPCELL_X1 PHY_54 ();
 AND2_X1 _08859_ (.A1(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_en ),
    .A2(clknet_3_5__leaf__00534_),
    .ZN(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ));
 AND2_X1 _08860_ (.A1(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_en ),
    .A2(clknet_3_0__leaf__00534_),
    .ZN(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ));
 AND2_X1 _08861_ (.A1(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_en ),
    .A2(clknet_3_3__leaf__00534_),
    .ZN(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ));
 AND2_X1 _08862_ (.A1(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_en ),
    .A2(clknet_3_1__leaf__00534_),
    .ZN(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ));
 AND2_X1 _08863_ (.A1(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_en ),
    .A2(clknet_3_1__leaf__00534_),
    .ZN(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ));
 AND2_X1 _08864_ (.A1(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_en ),
    .A2(clknet_3_3__leaf__00534_),
    .ZN(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ));
 AND2_X1 _08865_ (.A1(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_en ),
    .A2(clknet_3_4__leaf__00534_),
    .ZN(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ));
 AND2_X1 _08866_ (.A1(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_en ),
    .A2(clknet_3_3__leaf__00534_),
    .ZN(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ));
 AND2_X1 _08867_ (.A1(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_en ),
    .A2(clknet_3_1__leaf__00534_),
    .ZN(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ));
 TAPCELL_X1 PHY_53 ();
 AND2_X1 _08869_ (.A1(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_en ),
    .A2(clknet_3_6__leaf__00534_),
    .ZN(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ));
 AND2_X1 _08870_ (.A1(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_en ),
    .A2(clknet_3_4__leaf__00534_),
    .ZN(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ));
 AND2_X1 _08871_ (.A1(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_en ),
    .A2(clknet_3_7__leaf__00534_),
    .ZN(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ));
 AND2_X1 _08872_ (.A1(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_en ),
    .A2(clknet_3_2__leaf__00534_),
    .ZN(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ));
 AND2_X1 _08873_ (.A1(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_en ),
    .A2(clknet_3_0__leaf__00534_),
    .ZN(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ));
 AND2_X1 _08874_ (.A1(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_en ),
    .A2(clknet_3_2__leaf__00534_),
    .ZN(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ));
 AND2_X1 _08875_ (.A1(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_en ),
    .A2(clknet_3_2__leaf__00534_),
    .ZN(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ));
 AND2_X1 _08876_ (.A1(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_en ),
    .A2(clknet_3_0__leaf__00534_),
    .ZN(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ));
 AND2_X1 _08877_ (.A1(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_en ),
    .A2(clknet_3_6__leaf__00534_),
    .ZN(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ));
 AND2_X1 _08878_ (.A1(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_en ),
    .A2(clknet_3_2__leaf__00534_),
    .ZN(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ));
 TAPCELL_X1 PHY_52 ();
 AND2_X1 _08880_ (.A1(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_en ),
    .A2(clknet_3_2__leaf__00534_),
    .ZN(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ));
 AND2_X1 _08881_ (.A1(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_en ),
    .A2(clknet_3_3__leaf__00534_),
    .ZN(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ));
 AND2_X1 _08882_ (.A1(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_en ),
    .A2(clknet_3_7__leaf__00534_),
    .ZN(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ));
 AND2_X1 _08883_ (.A1(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_en ),
    .A2(clknet_3_2__leaf__00534_),
    .ZN(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ));
 AND2_X1 _08884_ (.A1(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_en ),
    .A2(clknet_3_4__leaf__00534_),
    .ZN(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ));
 AND2_X1 _08885_ (.A1(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_en ),
    .A2(clknet_3_1__leaf__00534_),
    .ZN(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ));
 AND2_X1 _08886_ (.A1(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_en ),
    .A2(clknet_3_5__leaf__00534_),
    .ZN(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ));
 AND2_X1 _08887_ (.A1(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_en ),
    .A2(clknet_3_1__leaf__00534_),
    .ZN(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ));
 AND2_X1 _08888_ (.A1(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_en ),
    .A2(clknet_3_4__leaf__00534_),
    .ZN(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ));
 AND2_X1 _08889_ (.A1(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_en ),
    .A2(clknet_3_7__leaf__00534_),
    .ZN(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ));
 AND2_X1 _08890_ (.A1(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_en ),
    .A2(clknet_3_6__leaf__00534_),
    .ZN(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ));
 AND2_X1 _08891_ (.A1(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_en ),
    .A2(clknet_3_6__leaf__00534_),
    .ZN(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ));
 AND2_X1 _08892_ (.A1(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_en ),
    .A2(clknet_3_4__leaf__00534_),
    .ZN(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ));
 AND2_X1 _08893_ (.A1(\lut.gen_sub_units_scm.__14.sub_unit_i.cg_we_global.clk_en ),
    .A2(clknet_2_1__leaf__00532_),
    .ZN(_00537_));
 TAPCELL_X1 PHY_51 ();
 AND2_X1 _08895_ (.A1(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_en ),
    .A2(clknet_3_6__leaf__00537_),
    .ZN(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ));
 AND2_X1 _08896_ (.A1(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_en ),
    .A2(clknet_3_2__leaf__00537_),
    .ZN(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ));
 AND2_X1 _08897_ (.A1(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_en ),
    .A2(clknet_3_0__leaf__00537_),
    .ZN(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ));
 AND2_X1 _08898_ (.A1(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_en ),
    .A2(clknet_3_0__leaf__00537_),
    .ZN(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ));
 AND2_X1 _08899_ (.A1(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_en ),
    .A2(clknet_3_7__leaf__00537_),
    .ZN(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ));
 AND2_X1 _08900_ (.A1(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_en ),
    .A2(clknet_3_4__leaf__00537_),
    .ZN(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ));
 AND2_X1 _08901_ (.A1(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_en ),
    .A2(clknet_3_2__leaf__00537_),
    .ZN(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ));
 AND2_X1 _08902_ (.A1(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_en ),
    .A2(clknet_3_1__leaf__00537_),
    .ZN(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ));
 AND2_X1 _08903_ (.A1(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_en ),
    .A2(clknet_3_2__leaf__00537_),
    .ZN(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ));
 TAPCELL_X1 PHY_50 ();
 AND2_X1 _08905_ (.A1(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_en ),
    .A2(clknet_3_5__leaf__00537_),
    .ZN(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ));
 AND2_X1 _08906_ (.A1(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_en ),
    .A2(clknet_3_5__leaf__00537_),
    .ZN(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ));
 AND2_X1 _08907_ (.A1(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_en ),
    .A2(clknet_3_2__leaf__00537_),
    .ZN(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ));
 AND2_X1 _08908_ (.A1(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_en ),
    .A2(clknet_3_6__leaf__00537_),
    .ZN(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ));
 AND2_X1 _08909_ (.A1(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_en ),
    .A2(clknet_3_4__leaf__00537_),
    .ZN(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ));
 AND2_X1 _08910_ (.A1(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_en ),
    .A2(clknet_3_5__leaf__00537_),
    .ZN(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ));
 AND2_X1 _08911_ (.A1(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_en ),
    .A2(clknet_3_4__leaf__00537_),
    .ZN(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ));
 AND2_X1 _08912_ (.A1(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_en ),
    .A2(clknet_3_5__leaf__00537_),
    .ZN(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ));
 AND2_X1 _08913_ (.A1(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_en ),
    .A2(clknet_3_0__leaf__00537_),
    .ZN(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ));
 AND2_X1 _08914_ (.A1(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_en ),
    .A2(clknet_3_3__leaf__00537_),
    .ZN(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ));
 TAPCELL_X1 PHY_49 ();
 AND2_X1 _08916_ (.A1(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_en ),
    .A2(clknet_3_1__leaf__00537_),
    .ZN(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ));
 AND2_X1 _08917_ (.A1(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_en ),
    .A2(clknet_3_6__leaf__00537_),
    .ZN(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ));
 AND2_X1 _08918_ (.A1(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_en ),
    .A2(clknet_3_4__leaf__00537_),
    .ZN(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ));
 AND2_X1 _08919_ (.A1(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_en ),
    .A2(clknet_3_5__leaf__00537_),
    .ZN(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ));
 AND2_X1 _08920_ (.A1(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_en ),
    .A2(clknet_3_7__leaf__00537_),
    .ZN(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ));
 AND2_X1 _08921_ (.A1(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_en ),
    .A2(clknet_3_1__leaf__00537_),
    .ZN(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ));
 AND2_X1 _08922_ (.A1(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_en ),
    .A2(clknet_3_1__leaf__00537_),
    .ZN(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ));
 AND2_X1 _08923_ (.A1(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_en ),
    .A2(clknet_3_5__leaf__00537_),
    .ZN(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ));
 AND2_X1 _08924_ (.A1(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_en ),
    .A2(clknet_3_1__leaf__00537_),
    .ZN(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ));
 AND2_X1 _08925_ (.A1(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_en ),
    .A2(clknet_3_3__leaf__00537_),
    .ZN(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ));
 AND2_X1 _08926_ (.A1(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_en ),
    .A2(clknet_3_7__leaf__00537_),
    .ZN(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ));
 AND2_X1 _08927_ (.A1(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_en ),
    .A2(clknet_3_7__leaf__00537_),
    .ZN(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ));
 AND2_X1 _08928_ (.A1(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_en ),
    .A2(clknet_3_0__leaf__00537_),
    .ZN(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ));
 AND2_X1 _08929_ (.A1(\lut.gen_sub_units_scm.__13.sub_unit_i.cg_we_global.clk_en ),
    .A2(clknet_2_3__leaf__00532_),
    .ZN(_00540_));
 TAPCELL_X1 PHY_48 ();
 AND2_X1 _08931_ (.A1(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_en ),
    .A2(clknet_3_4__leaf__00540_),
    .ZN(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ));
 AND2_X1 _08932_ (.A1(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_en ),
    .A2(clknet_3_6__leaf__00540_),
    .ZN(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ));
 AND2_X1 _08933_ (.A1(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_en ),
    .A2(clknet_3_2__leaf__00540_),
    .ZN(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ));
 AND2_X1 _08934_ (.A1(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_en ),
    .A2(clknet_3_5__leaf__00540_),
    .ZN(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ));
 AND2_X1 _08935_ (.A1(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_en ),
    .A2(clknet_3_3__leaf__00540_),
    .ZN(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ));
 AND2_X1 _08936_ (.A1(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_en ),
    .A2(clknet_3_2__leaf__00540_),
    .ZN(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ));
 AND2_X1 _08937_ (.A1(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_en ),
    .A2(clknet_3_2__leaf__00540_),
    .ZN(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ));
 AND2_X1 _08938_ (.A1(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_en ),
    .A2(clknet_3_1__leaf__00540_),
    .ZN(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ));
 AND2_X1 _08939_ (.A1(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_en ),
    .A2(clknet_3_6__leaf__00540_),
    .ZN(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ));
 TAPCELL_X1 PHY_47 ();
 AND2_X1 _08941_ (.A1(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_en ),
    .A2(clknet_3_3__leaf__00540_),
    .ZN(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ));
 AND2_X1 _08942_ (.A1(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_en ),
    .A2(clknet_3_7__leaf__00540_),
    .ZN(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ));
 AND2_X1 _08943_ (.A1(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_en ),
    .A2(clknet_3_3__leaf__00540_),
    .ZN(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ));
 AND2_X1 _08944_ (.A1(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_en ),
    .A2(clknet_3_1__leaf__00540_),
    .ZN(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ));
 AND2_X1 _08945_ (.A1(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_en ),
    .A2(clknet_3_2__leaf__00540_),
    .ZN(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ));
 AND2_X1 _08946_ (.A1(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_en ),
    .A2(clknet_3_4__leaf__00540_),
    .ZN(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ));
 AND2_X1 _08947_ (.A1(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_en ),
    .A2(clknet_3_0__leaf__00540_),
    .ZN(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ));
 AND2_X1 _08948_ (.A1(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_en ),
    .A2(clknet_3_7__leaf__00540_),
    .ZN(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ));
 AND2_X1 _08949_ (.A1(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_en ),
    .A2(clknet_3_5__leaf__00540_),
    .ZN(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ));
 AND2_X1 _08950_ (.A1(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_en ),
    .A2(clknet_3_6__leaf__00540_),
    .ZN(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ));
 TAPCELL_X1 PHY_46 ();
 AND2_X1 _08952_ (.A1(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_en ),
    .A2(clknet_3_3__leaf__00540_),
    .ZN(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ));
 AND2_X1 _08953_ (.A1(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_en ),
    .A2(clknet_3_0__leaf__00540_),
    .ZN(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ));
 AND2_X1 _08954_ (.A1(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_en ),
    .A2(clknet_3_0__leaf__00540_),
    .ZN(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ));
 AND2_X1 _08955_ (.A1(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_en ),
    .A2(clknet_3_3__leaf__00540_),
    .ZN(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ));
 AND2_X1 _08956_ (.A1(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_en ),
    .A2(clknet_3_7__leaf__00540_),
    .ZN(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ));
 AND2_X1 _08957_ (.A1(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_en ),
    .A2(clknet_3_2__leaf__00540_),
    .ZN(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ));
 AND2_X1 _08958_ (.A1(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_en ),
    .A2(clknet_3_0__leaf__00540_),
    .ZN(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ));
 AND2_X1 _08959_ (.A1(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_en ),
    .A2(clknet_3_2__leaf__00540_),
    .ZN(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ));
 AND2_X1 _08960_ (.A1(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_en ),
    .A2(clknet_3_1__leaf__00540_),
    .ZN(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ));
 AND2_X1 _08961_ (.A1(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_en ),
    .A2(clknet_3_5__leaf__00540_),
    .ZN(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ));
 AND2_X1 _08962_ (.A1(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_en ),
    .A2(clknet_3_7__leaf__00540_),
    .ZN(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ));
 AND2_X1 _08963_ (.A1(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_en ),
    .A2(clknet_3_1__leaf__00540_),
    .ZN(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ));
 AND2_X1 _08964_ (.A1(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_en ),
    .A2(clknet_3_7__leaf__00540_),
    .ZN(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ));
 AND2_X1 _08965_ (.A1(\lut.gen_sub_units_scm.__12.sub_unit_i.cg_we_global.clk_en ),
    .A2(clknet_2_1__leaf__00532_),
    .ZN(_00543_));
 TAPCELL_X1 PHY_45 ();
 AND2_X1 _08967_ (.A1(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_en ),
    .A2(clknet_3_5__leaf__00543_),
    .ZN(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ));
 AND2_X1 _08968_ (.A1(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_en ),
    .A2(clknet_3_7__leaf__00543_),
    .ZN(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ));
 AND2_X1 _08969_ (.A1(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_en ),
    .A2(clknet_3_4__leaf__00543_),
    .ZN(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ));
 AND2_X1 _08970_ (.A1(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_en ),
    .A2(clknet_3_7__leaf__00543_),
    .ZN(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ));
 AND2_X1 _08971_ (.A1(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_en ),
    .A2(clknet_3_2__leaf__00543_),
    .ZN(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ));
 AND2_X1 _08972_ (.A1(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_en ),
    .A2(clknet_3_0__leaf__00543_),
    .ZN(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ));
 AND2_X1 _08973_ (.A1(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_en ),
    .A2(clknet_3_3__leaf__00543_),
    .ZN(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ));
 AND2_X1 _08974_ (.A1(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_en ),
    .A2(clknet_3_3__leaf__00543_),
    .ZN(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ));
 AND2_X1 _08975_ (.A1(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_en ),
    .A2(clknet_3_2__leaf__00543_),
    .ZN(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ));
 TAPCELL_X1 PHY_44 ();
 AND2_X1 _08977_ (.A1(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_en ),
    .A2(clknet_3_3__leaf__00543_),
    .ZN(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ));
 AND2_X1 _08978_ (.A1(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_en ),
    .A2(clknet_3_6__leaf__00543_),
    .ZN(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ));
 AND2_X1 _08979_ (.A1(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_en ),
    .A2(clknet_3_1__leaf__00543_),
    .ZN(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ));
 AND2_X1 _08980_ (.A1(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_en ),
    .A2(clknet_3_4__leaf__00543_),
    .ZN(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ));
 AND2_X1 _08981_ (.A1(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_en ),
    .A2(clknet_3_2__leaf__00543_),
    .ZN(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ));
 AND2_X1 _08982_ (.A1(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_en ),
    .A2(clknet_3_5__leaf__00543_),
    .ZN(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ));
 AND2_X1 _08983_ (.A1(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_en ),
    .A2(clknet_3_3__leaf__00543_),
    .ZN(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ));
 AND2_X1 _08984_ (.A1(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_en ),
    .A2(clknet_3_7__leaf__00543_),
    .ZN(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ));
 AND2_X1 _08985_ (.A1(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_en ),
    .A2(clknet_3_4__leaf__00543_),
    .ZN(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ));
 AND2_X1 _08986_ (.A1(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_en ),
    .A2(clknet_3_7__leaf__00543_),
    .ZN(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ));
 TAPCELL_X1 PHY_43 ();
 AND2_X1 _08988_ (.A1(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_en ),
    .A2(clknet_3_6__leaf__00543_),
    .ZN(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ));
 AND2_X1 _08989_ (.A1(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_en ),
    .A2(clknet_3_6__leaf__00543_),
    .ZN(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ));
 AND2_X1 _08990_ (.A1(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_en ),
    .A2(clknet_3_1__leaf__00543_),
    .ZN(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ));
 AND2_X1 _08991_ (.A1(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_en ),
    .A2(clknet_3_7__leaf__00543_),
    .ZN(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ));
 AND2_X1 _08992_ (.A1(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_en ),
    .A2(clknet_3_1__leaf__00543_),
    .ZN(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ));
 AND2_X1 _08993_ (.A1(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_en ),
    .A2(clknet_3_4__leaf__00543_),
    .ZN(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ));
 AND2_X1 _08994_ (.A1(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_en ),
    .A2(clknet_3_0__leaf__00543_),
    .ZN(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ));
 AND2_X1 _08995_ (.A1(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_en ),
    .A2(clknet_3_1__leaf__00543_),
    .ZN(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ));
 AND2_X1 _08996_ (.A1(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_en ),
    .A2(clknet_3_3__leaf__00543_),
    .ZN(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ));
 AND2_X1 _08997_ (.A1(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_en ),
    .A2(clknet_3_2__leaf__00543_),
    .ZN(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ));
 AND2_X1 _08998_ (.A1(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_en ),
    .A2(clknet_3_1__leaf__00543_),
    .ZN(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ));
 AND2_X1 _08999_ (.A1(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_en ),
    .A2(clknet_3_0__leaf__00543_),
    .ZN(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ));
 AND2_X1 _09000_ (.A1(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_en ),
    .A2(clknet_3_2__leaf__00543_),
    .ZN(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ));
 AND2_X1 _09001_ (.A1(\lut.gen_sub_units_scm.__11.sub_unit_i.cg_we_global.clk_en ),
    .A2(clknet_2_3__leaf__00532_),
    .ZN(_00546_));
 TAPCELL_X1 PHY_42 ();
 AND2_X1 _09003_ (.A1(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_en ),
    .A2(clknet_3_4__leaf__00546_),
    .ZN(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ));
 AND2_X1 _09004_ (.A1(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_en ),
    .A2(clknet_3_3__leaf__00546_),
    .ZN(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ));
 AND2_X1 _09005_ (.A1(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_en ),
    .A2(clknet_3_2__leaf__00546_),
    .ZN(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ));
 AND2_X1 _09006_ (.A1(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_en ),
    .A2(clknet_3_6__leaf__00546_),
    .ZN(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ));
 AND2_X1 _09007_ (.A1(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_en ),
    .A2(clknet_3_4__leaf__00546_),
    .ZN(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ));
 AND2_X1 _09008_ (.A1(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_en ),
    .A2(clknet_3_7__leaf__00546_),
    .ZN(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ));
 AND2_X1 _09009_ (.A1(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_en ),
    .A2(clknet_3_0__leaf__00546_),
    .ZN(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ));
 AND2_X1 _09010_ (.A1(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_en ),
    .A2(clknet_3_7__leaf__00546_),
    .ZN(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ));
 AND2_X1 _09011_ (.A1(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_en ),
    .A2(clknet_3_3__leaf__00546_),
    .ZN(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ));
 TAPCELL_X1 PHY_41 ();
 AND2_X1 _09013_ (.A1(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_en ),
    .A2(clknet_3_5__leaf__00546_),
    .ZN(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ));
 AND2_X1 _09014_ (.A1(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_en ),
    .A2(clknet_3_6__leaf__00546_),
    .ZN(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ));
 AND2_X1 _09015_ (.A1(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_en ),
    .A2(clknet_3_2__leaf__00546_),
    .ZN(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ));
 AND2_X1 _09016_ (.A1(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_en ),
    .A2(clknet_3_2__leaf__00546_),
    .ZN(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ));
 AND2_X1 _09017_ (.A1(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_en ),
    .A2(clknet_3_4__leaf__00546_),
    .ZN(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ));
 AND2_X1 _09018_ (.A1(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_en ),
    .A2(clknet_3_2__leaf__00546_),
    .ZN(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ));
 AND2_X1 _09019_ (.A1(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_en ),
    .A2(clknet_3_0__leaf__00546_),
    .ZN(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ));
 AND2_X1 _09020_ (.A1(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_en ),
    .A2(clknet_3_0__leaf__00546_),
    .ZN(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ));
 AND2_X1 _09021_ (.A1(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_en ),
    .A2(clknet_3_6__leaf__00546_),
    .ZN(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ));
 AND2_X1 _09022_ (.A1(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_en ),
    .A2(clknet_3_3__leaf__00546_),
    .ZN(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ));
 TAPCELL_X1 PHY_40 ();
 AND2_X1 _09024_ (.A1(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_en ),
    .A2(clknet_3_1__leaf__00546_),
    .ZN(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ));
 AND2_X1 _09025_ (.A1(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_en ),
    .A2(clknet_3_7__leaf__00546_),
    .ZN(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ));
 AND2_X1 _09026_ (.A1(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_en ),
    .A2(clknet_3_5__leaf__00546_),
    .ZN(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ));
 AND2_X1 _09027_ (.A1(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_en ),
    .A2(clknet_3_2__leaf__00546_),
    .ZN(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ));
 AND2_X1 _09028_ (.A1(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_en ),
    .A2(clknet_3_3__leaf__00546_),
    .ZN(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ));
 AND2_X1 _09029_ (.A1(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_en ),
    .A2(clknet_3_3__leaf__00546_),
    .ZN(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ));
 AND2_X1 _09030_ (.A1(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_en ),
    .A2(clknet_3_5__leaf__00546_),
    .ZN(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ));
 AND2_X1 _09031_ (.A1(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_en ),
    .A2(clknet_3_6__leaf__00546_),
    .ZN(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ));
 AND2_X1 _09032_ (.A1(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_en ),
    .A2(clknet_3_4__leaf__00546_),
    .ZN(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ));
 AND2_X1 _09033_ (.A1(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_en ),
    .A2(clknet_3_0__leaf__00546_),
    .ZN(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ));
 AND2_X1 _09034_ (.A1(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_en ),
    .A2(clknet_3_0__leaf__00546_),
    .ZN(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ));
 AND2_X1 _09035_ (.A1(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_en ),
    .A2(clknet_3_2__leaf__00546_),
    .ZN(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ));
 AND2_X1 _09036_ (.A1(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_en ),
    .A2(clknet_3_3__leaf__00546_),
    .ZN(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ));
 AND2_X1 _09037_ (.A1(\lut.gen_sub_units_scm.__10.sub_unit_i.cg_we_global.clk_en ),
    .A2(clknet_2_0__leaf__00532_),
    .ZN(_00549_));
 TAPCELL_X1 PHY_39 ();
 AND2_X1 _09039_ (.A1(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_en ),
    .A2(clknet_3_7__leaf__00549_),
    .ZN(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ));
 AND2_X1 _09040_ (.A1(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_en ),
    .A2(clknet_3_1__leaf__00549_),
    .ZN(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ));
 AND2_X1 _09041_ (.A1(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_en ),
    .A2(clknet_3_0__leaf__00549_),
    .ZN(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ));
 AND2_X1 _09042_ (.A1(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_en ),
    .A2(clknet_3_1__leaf__00549_),
    .ZN(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ));
 AND2_X1 _09043_ (.A1(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_en ),
    .A2(clknet_3_0__leaf__00549_),
    .ZN(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ));
 AND2_X1 _09044_ (.A1(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_en ),
    .A2(clknet_3_4__leaf__00549_),
    .ZN(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ));
 AND2_X1 _09045_ (.A1(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_en ),
    .A2(clknet_3_3__leaf__00549_),
    .ZN(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ));
 AND2_X1 _09046_ (.A1(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_en ),
    .A2(clknet_3_0__leaf__00549_),
    .ZN(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ));
 AND2_X1 _09047_ (.A1(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_en ),
    .A2(clknet_3_6__leaf__00549_),
    .ZN(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ));
 TAPCELL_X1 PHY_38 ();
 AND2_X1 _09049_ (.A1(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_en ),
    .A2(clknet_3_4__leaf__00549_),
    .ZN(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ));
 AND2_X1 _09050_ (.A1(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_en ),
    .A2(clknet_3_2__leaf__00549_),
    .ZN(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ));
 AND2_X1 _09051_ (.A1(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_en ),
    .A2(clknet_3_2__leaf__00549_),
    .ZN(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ));
 AND2_X1 _09052_ (.A1(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_en ),
    .A2(clknet_3_1__leaf__00549_),
    .ZN(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ));
 AND2_X1 _09053_ (.A1(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_en ),
    .A2(clknet_3_5__leaf__00549_),
    .ZN(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ));
 AND2_X1 _09054_ (.A1(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_en ),
    .A2(clknet_3_4__leaf__00549_),
    .ZN(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ));
 AND2_X1 _09055_ (.A1(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_en ),
    .A2(clknet_3_1__leaf__00549_),
    .ZN(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ));
 AND2_X1 _09056_ (.A1(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_en ),
    .A2(clknet_3_5__leaf__00549_),
    .ZN(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ));
 AND2_X1 _09057_ (.A1(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_en ),
    .A2(clknet_3_2__leaf__00549_),
    .ZN(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ));
 AND2_X1 _09058_ (.A1(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_en ),
    .A2(clknet_3_5__leaf__00549_),
    .ZN(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ));
 TAPCELL_X1 PHY_37 ();
 AND2_X1 _09060_ (.A1(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_en ),
    .A2(clknet_3_1__leaf__00549_),
    .ZN(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ));
 AND2_X1 _09061_ (.A1(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_en ),
    .A2(clknet_3_5__leaf__00549_),
    .ZN(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ));
 AND2_X1 _09062_ (.A1(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_en ),
    .A2(clknet_3_3__leaf__00549_),
    .ZN(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ));
 AND2_X1 _09063_ (.A1(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_en ),
    .A2(clknet_3_7__leaf__00549_),
    .ZN(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ));
 AND2_X1 _09064_ (.A1(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_en ),
    .A2(clknet_3_3__leaf__00549_),
    .ZN(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ));
 AND2_X1 _09065_ (.A1(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_en ),
    .A2(clknet_3_4__leaf__00549_),
    .ZN(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ));
 AND2_X1 _09066_ (.A1(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_en ),
    .A2(clknet_3_3__leaf__00549_),
    .ZN(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ));
 AND2_X1 _09067_ (.A1(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_en ),
    .A2(clknet_3_1__leaf__00549_),
    .ZN(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ));
 AND2_X1 _09068_ (.A1(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_en ),
    .A2(clknet_3_7__leaf__00549_),
    .ZN(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ));
 AND2_X1 _09069_ (.A1(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_en ),
    .A2(clknet_3_6__leaf__00549_),
    .ZN(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ));
 AND2_X1 _09070_ (.A1(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_en ),
    .A2(clknet_3_0__leaf__00549_),
    .ZN(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ));
 AND2_X1 _09071_ (.A1(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_en ),
    .A2(clknet_3_3__leaf__00549_),
    .ZN(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ));
 AND2_X1 _09072_ (.A1(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_en ),
    .A2(clknet_3_0__leaf__00549_),
    .ZN(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ));
 AND2_X1 _09073_ (.A1(\lut.gen_sub_units_scm.__9.sub_unit_i.cg_we_global.clk_en ),
    .A2(clknet_2_1__leaf__00532_),
    .ZN(_00552_));
 TAPCELL_X1 PHY_36 ();
 AND2_X1 _09075_ (.A1(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_en ),
    .A2(clknet_3_6__leaf__00552_),
    .ZN(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ));
 AND2_X1 _09076_ (.A1(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_en ),
    .A2(clknet_3_2__leaf__00552_),
    .ZN(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ));
 AND2_X1 _09077_ (.A1(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_en ),
    .A2(clknet_3_7__leaf__00552_),
    .ZN(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ));
 AND2_X1 _09078_ (.A1(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_en ),
    .A2(clknet_3_2__leaf__00552_),
    .ZN(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ));
 AND2_X1 _09079_ (.A1(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_en ),
    .A2(clknet_3_0__leaf__00552_),
    .ZN(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ));
 AND2_X1 _09080_ (.A1(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_en ),
    .A2(clknet_3_3__leaf__00552_),
    .ZN(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ));
 AND2_X1 _09081_ (.A1(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_en ),
    .A2(clknet_3_5__leaf__00552_),
    .ZN(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ));
 AND2_X1 _09082_ (.A1(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_en ),
    .A2(clknet_3_2__leaf__00552_),
    .ZN(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ));
 AND2_X1 _09083_ (.A1(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_en ),
    .A2(clknet_3_0__leaf__00552_),
    .ZN(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ));
 TAPCELL_X1 PHY_35 ();
 AND2_X1 _09085_ (.A1(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_en ),
    .A2(clknet_3_5__leaf__00552_),
    .ZN(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ));
 AND2_X1 _09086_ (.A1(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_en ),
    .A2(clknet_3_0__leaf__00552_),
    .ZN(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ));
 AND2_X1 _09087_ (.A1(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_en ),
    .A2(clknet_3_7__leaf__00552_),
    .ZN(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ));
 AND2_X1 _09088_ (.A1(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_en ),
    .A2(clknet_3_7__leaf__00552_),
    .ZN(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ));
 AND2_X1 _09089_ (.A1(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_en ),
    .A2(clknet_3_4__leaf__00552_),
    .ZN(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ));
 AND2_X1 _09090_ (.A1(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_en ),
    .A2(clknet_3_6__leaf__00552_),
    .ZN(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ));
 AND2_X1 _09091_ (.A1(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_en ),
    .A2(clknet_3_1__leaf__00552_),
    .ZN(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ));
 AND2_X1 _09092_ (.A1(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_en ),
    .A2(clknet_3_1__leaf__00552_),
    .ZN(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ));
 AND2_X1 _09093_ (.A1(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_en ),
    .A2(clknet_3_6__leaf__00552_),
    .ZN(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ));
 AND2_X1 _09094_ (.A1(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_en ),
    .A2(clknet_3_7__leaf__00552_),
    .ZN(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ));
 TAPCELL_X1 PHY_34 ();
 AND2_X1 _09096_ (.A1(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_en ),
    .A2(clknet_3_4__leaf__00552_),
    .ZN(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ));
 AND2_X1 _09097_ (.A1(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_en ),
    .A2(clknet_3_4__leaf__00552_),
    .ZN(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ));
 AND2_X1 _09098_ (.A1(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_en ),
    .A2(clknet_3_7__leaf__00552_),
    .ZN(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ));
 AND2_X1 _09099_ (.A1(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_en ),
    .A2(clknet_3_5__leaf__00552_),
    .ZN(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ));
 AND2_X1 _09100_ (.A1(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_en ),
    .A2(clknet_3_1__leaf__00552_),
    .ZN(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ));
 AND2_X1 _09101_ (.A1(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_en ),
    .A2(clknet_3_3__leaf__00552_),
    .ZN(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ));
 AND2_X1 _09102_ (.A1(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_en ),
    .A2(clknet_3_5__leaf__00552_),
    .ZN(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ));
 AND2_X1 _09103_ (.A1(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_en ),
    .A2(clknet_3_5__leaf__00552_),
    .ZN(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ));
 AND2_X1 _09104_ (.A1(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_en ),
    .A2(clknet_3_3__leaf__00552_),
    .ZN(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ));
 AND2_X1 _09105_ (.A1(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_en ),
    .A2(clknet_3_6__leaf__00552_),
    .ZN(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ));
 AND2_X1 _09106_ (.A1(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_en ),
    .A2(clknet_3_1__leaf__00552_),
    .ZN(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ));
 AND2_X1 _09107_ (.A1(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_en ),
    .A2(clknet_3_4__leaf__00552_),
    .ZN(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ));
 AND2_X1 _09108_ (.A1(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_en ),
    .A2(clknet_3_0__leaf__00552_),
    .ZN(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ));
 AND2_X1 _09109_ (.A1(\lut.gen_sub_units_scm.__8.sub_unit_i.cg_we_global.clk_en ),
    .A2(clknet_2_0__leaf__00532_),
    .ZN(_00555_));
 TAPCELL_X1 PHY_33 ();
 AND2_X1 _09111_ (.A1(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_en ),
    .A2(clknet_3_7__leaf__00555_),
    .ZN(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ));
 AND2_X1 _09112_ (.A1(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_en ),
    .A2(clknet_3_0__leaf__00555_),
    .ZN(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ));
 AND2_X1 _09113_ (.A1(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_en ),
    .A2(clknet_3_3__leaf__00555_),
    .ZN(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ));
 AND2_X1 _09114_ (.A1(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_en ),
    .A2(clknet_3_7__leaf__00555_),
    .ZN(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ));
 AND2_X1 _09115_ (.A1(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_en ),
    .A2(clknet_3_1__leaf__00555_),
    .ZN(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ));
 AND2_X1 _09116_ (.A1(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_en ),
    .A2(clknet_3_1__leaf__00555_),
    .ZN(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ));
 AND2_X1 _09117_ (.A1(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_en ),
    .A2(clknet_3_4__leaf__00555_),
    .ZN(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ));
 AND2_X1 _09118_ (.A1(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_en ),
    .A2(clknet_3_3__leaf__00555_),
    .ZN(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ));
 AND2_X1 _09119_ (.A1(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_en ),
    .A2(clknet_3_1__leaf__00555_),
    .ZN(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ));
 TAPCELL_X1 PHY_32 ();
 AND2_X1 _09121_ (.A1(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_en ),
    .A2(clknet_3_4__leaf__00555_),
    .ZN(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ));
 AND2_X1 _09122_ (.A1(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_en ),
    .A2(clknet_3_4__leaf__00555_),
    .ZN(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ));
 AND2_X1 _09123_ (.A1(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_en ),
    .A2(clknet_3_6__leaf__00555_),
    .ZN(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ));
 AND2_X1 _09124_ (.A1(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_en ),
    .A2(clknet_3_3__leaf__00555_),
    .ZN(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ));
 AND2_X1 _09125_ (.A1(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_en ),
    .A2(clknet_3_0__leaf__00555_),
    .ZN(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ));
 AND2_X1 _09126_ (.A1(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_en ),
    .A2(clknet_3_2__leaf__00555_),
    .ZN(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ));
 AND2_X1 _09127_ (.A1(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_en ),
    .A2(clknet_3_2__leaf__00555_),
    .ZN(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ));
 AND2_X1 _09128_ (.A1(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_en ),
    .A2(clknet_3_2__leaf__00555_),
    .ZN(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ));
 AND2_X1 _09129_ (.A1(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_en ),
    .A2(clknet_3_6__leaf__00555_),
    .ZN(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ));
 AND2_X1 _09130_ (.A1(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_en ),
    .A2(clknet_3_2__leaf__00555_),
    .ZN(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ));
 TAPCELL_X1 PHY_31 ();
 AND2_X1 _09132_ (.A1(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_en ),
    .A2(clknet_3_0__leaf__00555_),
    .ZN(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ));
 AND2_X1 _09133_ (.A1(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_en ),
    .A2(clknet_3_1__leaf__00555_),
    .ZN(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ));
 AND2_X1 _09134_ (.A1(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_en ),
    .A2(clknet_3_7__leaf__00555_),
    .ZN(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ));
 AND2_X1 _09135_ (.A1(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_en ),
    .A2(clknet_3_2__leaf__00555_),
    .ZN(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ));
 AND2_X1 _09136_ (.A1(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_en ),
    .A2(clknet_3_1__leaf__00555_),
    .ZN(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ));
 AND2_X1 _09137_ (.A1(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_en ),
    .A2(clknet_3_3__leaf__00555_),
    .ZN(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ));
 AND2_X1 _09138_ (.A1(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_en ),
    .A2(clknet_3_5__leaf__00555_),
    .ZN(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ));
 AND2_X1 _09139_ (.A1(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_en ),
    .A2(clknet_3_0__leaf__00555_),
    .ZN(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ));
 AND2_X1 _09140_ (.A1(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_en ),
    .A2(clknet_3_5__leaf__00555_),
    .ZN(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ));
 AND2_X1 _09141_ (.A1(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_en ),
    .A2(clknet_3_4__leaf__00555_),
    .ZN(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ));
 AND2_X1 _09142_ (.A1(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_en ),
    .A2(clknet_3_3__leaf__00555_),
    .ZN(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ));
 AND2_X1 _09143_ (.A1(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_en ),
    .A2(clknet_3_4__leaf__00555_),
    .ZN(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ));
 AND2_X1 _09144_ (.A1(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_en ),
    .A2(clknet_3_5__leaf__00555_),
    .ZN(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ));
 AND2_X1 _09145_ (.A1(\lut.gen_sub_units_scm.__7.sub_unit_i.cg_we_global.clk_en ),
    .A2(clknet_2_0__leaf__00532_),
    .ZN(_00558_));
 TAPCELL_X1 PHY_30 ();
 AND2_X1 _09147_ (.A1(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_en ),
    .A2(clknet_3_5__leaf__00558_),
    .ZN(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ));
 AND2_X1 _09148_ (.A1(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_en ),
    .A2(clknet_3_3__leaf__00558_),
    .ZN(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ));
 AND2_X1 _09149_ (.A1(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_en ),
    .A2(clknet_3_0__leaf__00558_),
    .ZN(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ));
 AND2_X1 _09150_ (.A1(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_en ),
    .A2(clknet_3_6__leaf__00558_),
    .ZN(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ));
 AND2_X1 _09151_ (.A1(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_en ),
    .A2(clknet_3_1__leaf__00558_),
    .ZN(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ));
 AND2_X1 _09152_ (.A1(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_en ),
    .A2(clknet_3_5__leaf__00558_),
    .ZN(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ));
 AND2_X1 _09153_ (.A1(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_en ),
    .A2(clknet_3_6__leaf__00558_),
    .ZN(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ));
 AND2_X1 _09154_ (.A1(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_en ),
    .A2(clknet_3_0__leaf__00558_),
    .ZN(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ));
 AND2_X1 _09155_ (.A1(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_en ),
    .A2(clknet_3_2__leaf__00558_),
    .ZN(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ));
 TAPCELL_X1 PHY_29 ();
 AND2_X1 _09157_ (.A1(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_en ),
    .A2(clknet_3_6__leaf__00558_),
    .ZN(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ));
 AND2_X1 _09158_ (.A1(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_en ),
    .A2(clknet_3_5__leaf__00558_),
    .ZN(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ));
 AND2_X1 _09159_ (.A1(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_en ),
    .A2(clknet_3_4__leaf__00558_),
    .ZN(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ));
 AND2_X1 _09160_ (.A1(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_en ),
    .A2(clknet_3_0__leaf__00558_),
    .ZN(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ));
 AND2_X1 _09161_ (.A1(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_en ),
    .A2(clknet_3_7__leaf__00558_),
    .ZN(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ));
 AND2_X1 _09162_ (.A1(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_en ),
    .A2(clknet_3_3__leaf__00558_),
    .ZN(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ));
 AND2_X1 _09163_ (.A1(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_en ),
    .A2(clknet_3_6__leaf__00558_),
    .ZN(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ));
 AND2_X1 _09164_ (.A1(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_en ),
    .A2(clknet_3_5__leaf__00558_),
    .ZN(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ));
 AND2_X1 _09165_ (.A1(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_en ),
    .A2(clknet_3_4__leaf__00558_),
    .ZN(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ));
 AND2_X1 _09166_ (.A1(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_en ),
    .A2(clknet_3_2__leaf__00558_),
    .ZN(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ));
 TAPCELL_X1 PHY_28 ();
 AND2_X1 _09168_ (.A1(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_en ),
    .A2(clknet_3_3__leaf__00558_),
    .ZN(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ));
 AND2_X1 _09169_ (.A1(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_en ),
    .A2(clknet_3_2__leaf__00558_),
    .ZN(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ));
 AND2_X1 _09170_ (.A1(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_en ),
    .A2(clknet_3_4__leaf__00558_),
    .ZN(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ));
 AND2_X1 _09171_ (.A1(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_en ),
    .A2(clknet_3_4__leaf__00558_),
    .ZN(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ));
 AND2_X1 _09172_ (.A1(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_en ),
    .A2(clknet_3_2__leaf__00558_),
    .ZN(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ));
 AND2_X1 _09173_ (.A1(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_en ),
    .A2(clknet_3_1__leaf__00558_),
    .ZN(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ));
 AND2_X1 _09174_ (.A1(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_en ),
    .A2(clknet_3_5__leaf__00558_),
    .ZN(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ));
 AND2_X1 _09175_ (.A1(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_en ),
    .A2(clknet_3_2__leaf__00558_),
    .ZN(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ));
 AND2_X1 _09176_ (.A1(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_en ),
    .A2(clknet_3_2__leaf__00558_),
    .ZN(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ));
 AND2_X1 _09177_ (.A1(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_en ),
    .A2(clknet_3_7__leaf__00558_),
    .ZN(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ));
 AND2_X1 _09178_ (.A1(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_en ),
    .A2(clknet_3_7__leaf__00558_),
    .ZN(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ));
 AND2_X1 _09179_ (.A1(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_en ),
    .A2(clknet_3_0__leaf__00558_),
    .ZN(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ));
 AND2_X1 _09180_ (.A1(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_en ),
    .A2(clknet_3_4__leaf__00558_),
    .ZN(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ));
 AND2_X1 _09181_ (.A1(\lut.gen_sub_units_scm.__6.sub_unit_i.cg_we_global.clk_en ),
    .A2(clknet_2_0__leaf__00532_),
    .ZN(_00561_));
 TAPCELL_X1 PHY_27 ();
 AND2_X1 _09183_ (.A1(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_en ),
    .A2(clknet_3_3__leaf__00561_),
    .ZN(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ));
 AND2_X1 _09184_ (.A1(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_en ),
    .A2(clknet_3_1__leaf__00561_),
    .ZN(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ));
 AND2_X1 _09185_ (.A1(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_en ),
    .A2(clknet_3_3__leaf__00561_),
    .ZN(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ));
 AND2_X1 _09186_ (.A1(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_en ),
    .A2(clknet_3_4__leaf__00561_),
    .ZN(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ));
 AND2_X1 _09187_ (.A1(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_en ),
    .A2(clknet_3_2__leaf__00561_),
    .ZN(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ));
 AND2_X1 _09188_ (.A1(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_en ),
    .A2(clknet_3_1__leaf__00561_),
    .ZN(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ));
 AND2_X1 _09189_ (.A1(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_en ),
    .A2(clknet_3_7__leaf__00561_),
    .ZN(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ));
 AND2_X1 _09190_ (.A1(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_en ),
    .A2(clknet_3_6__leaf__00561_),
    .ZN(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ));
 AND2_X1 _09191_ (.A1(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_en ),
    .A2(clknet_3_2__leaf__00561_),
    .ZN(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ));
 TAPCELL_X1 PHY_26 ();
 AND2_X1 _09193_ (.A1(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_en ),
    .A2(clknet_3_2__leaf__00561_),
    .ZN(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ));
 AND2_X1 _09194_ (.A1(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_en ),
    .A2(clknet_3_0__leaf__00561_),
    .ZN(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ));
 AND2_X1 _09195_ (.A1(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_en ),
    .A2(clknet_3_7__leaf__00561_),
    .ZN(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ));
 AND2_X1 _09196_ (.A1(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_en ),
    .A2(clknet_3_6__leaf__00561_),
    .ZN(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ));
 AND2_X1 _09197_ (.A1(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_en ),
    .A2(clknet_3_1__leaf__00561_),
    .ZN(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ));
 AND2_X1 _09198_ (.A1(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_en ),
    .A2(clknet_3_7__leaf__00561_),
    .ZN(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ));
 AND2_X1 _09199_ (.A1(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_en ),
    .A2(clknet_3_5__leaf__00561_),
    .ZN(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ));
 AND2_X1 _09200_ (.A1(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_en ),
    .A2(clknet_3_5__leaf__00561_),
    .ZN(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ));
 AND2_X1 _09201_ (.A1(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_en ),
    .A2(clknet_3_5__leaf__00561_),
    .ZN(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ));
 AND2_X1 _09202_ (.A1(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_en ),
    .A2(clknet_3_1__leaf__00561_),
    .ZN(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ));
 TAPCELL_X1 PHY_25 ();
 AND2_X1 _09204_ (.A1(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_en ),
    .A2(clknet_3_0__leaf__00561_),
    .ZN(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ));
 AND2_X1 _09205_ (.A1(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_en ),
    .A2(clknet_3_5__leaf__00561_),
    .ZN(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ));
 AND2_X1 _09206_ (.A1(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_en ),
    .A2(clknet_3_5__leaf__00561_),
    .ZN(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ));
 AND2_X1 _09207_ (.A1(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_en ),
    .A2(clknet_3_1__leaf__00561_),
    .ZN(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ));
 AND2_X1 _09208_ (.A1(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_en ),
    .A2(clknet_3_5__leaf__00561_),
    .ZN(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ));
 AND2_X1 _09209_ (.A1(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_en ),
    .A2(clknet_3_6__leaf__00561_),
    .ZN(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ));
 AND2_X1 _09210_ (.A1(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_en ),
    .A2(clknet_3_0__leaf__00561_),
    .ZN(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ));
 AND2_X1 _09211_ (.A1(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_en ),
    .A2(clknet_3_0__leaf__00561_),
    .ZN(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ));
 AND2_X1 _09212_ (.A1(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_en ),
    .A2(clknet_3_7__leaf__00561_),
    .ZN(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ));
 AND2_X1 _09213_ (.A1(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_en ),
    .A2(clknet_3_2__leaf__00561_),
    .ZN(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ));
 AND2_X1 _09214_ (.A1(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_en ),
    .A2(clknet_3_1__leaf__00561_),
    .ZN(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ));
 AND2_X1 _09215_ (.A1(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_en ),
    .A2(clknet_3_2__leaf__00561_),
    .ZN(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ));
 AND2_X1 _09216_ (.A1(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_en ),
    .A2(clknet_3_0__leaf__00561_),
    .ZN(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ));
 AND2_X1 _09217_ (.A1(\lut.gen_sub_units_scm.__5.sub_unit_i.cg_we_global.clk_en ),
    .A2(clknet_2_2__leaf__00532_),
    .ZN(_00564_));
 TAPCELL_X1 PHY_24 ();
 AND2_X1 _09219_ (.A1(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_en ),
    .A2(clknet_3_1__leaf__00564_),
    .ZN(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ));
 AND2_X1 _09220_ (.A1(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_en ),
    .A2(clknet_3_6__leaf__00564_),
    .ZN(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ));
 AND2_X1 _09221_ (.A1(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_en ),
    .A2(clknet_3_3__leaf__00564_),
    .ZN(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ));
 AND2_X1 _09222_ (.A1(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_en ),
    .A2(clknet_3_1__leaf__00564_),
    .ZN(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ));
 AND2_X1 _09223_ (.A1(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_en ),
    .A2(clknet_3_2__leaf__00564_),
    .ZN(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ));
 AND2_X1 _09224_ (.A1(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_en ),
    .A2(clknet_3_2__leaf__00564_),
    .ZN(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ));
 AND2_X1 _09225_ (.A1(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_en ),
    .A2(clknet_3_5__leaf__00564_),
    .ZN(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ));
 AND2_X1 _09226_ (.A1(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_en ),
    .A2(clknet_3_7__leaf__00564_),
    .ZN(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ));
 AND2_X1 _09227_ (.A1(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_en ),
    .A2(clknet_3_1__leaf__00564_),
    .ZN(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ));
 TAPCELL_X1 PHY_23 ();
 AND2_X1 _09229_ (.A1(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_en ),
    .A2(clknet_3_3__leaf__00564_),
    .ZN(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ));
 AND2_X1 _09230_ (.A1(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_en ),
    .A2(clknet_3_4__leaf__00564_),
    .ZN(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ));
 AND2_X1 _09231_ (.A1(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_en ),
    .A2(clknet_3_3__leaf__00564_),
    .ZN(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ));
 AND2_X1 _09232_ (.A1(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_en ),
    .A2(clknet_3_3__leaf__00564_),
    .ZN(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ));
 AND2_X1 _09233_ (.A1(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_en ),
    .A2(clknet_3_0__leaf__00564_),
    .ZN(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ));
 AND2_X1 _09234_ (.A1(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_en ),
    .A2(clknet_3_3__leaf__00564_),
    .ZN(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ));
 AND2_X1 _09235_ (.A1(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_en ),
    .A2(clknet_3_3__leaf__00564_),
    .ZN(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ));
 AND2_X1 _09236_ (.A1(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_en ),
    .A2(clknet_3_4__leaf__00564_),
    .ZN(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ));
 AND2_X1 _09237_ (.A1(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_en ),
    .A2(clknet_3_3__leaf__00564_),
    .ZN(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ));
 AND2_X1 _09238_ (.A1(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_en ),
    .A2(clknet_3_0__leaf__00564_),
    .ZN(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ));
 TAPCELL_X1 PHY_22 ();
 AND2_X1 _09240_ (.A1(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_en ),
    .A2(clknet_3_7__leaf__00564_),
    .ZN(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ));
 AND2_X1 _09241_ (.A1(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_en ),
    .A2(clknet_3_7__leaf__00564_),
    .ZN(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ));
 AND2_X1 _09242_ (.A1(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_en ),
    .A2(clknet_3_2__leaf__00564_),
    .ZN(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ));
 AND2_X1 _09243_ (.A1(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_en ),
    .A2(clknet_3_0__leaf__00564_),
    .ZN(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ));
 AND2_X1 _09244_ (.A1(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_en ),
    .A2(clknet_3_7__leaf__00564_),
    .ZN(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ));
 AND2_X1 _09245_ (.A1(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_en ),
    .A2(clknet_3_5__leaf__00564_),
    .ZN(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ));
 AND2_X1 _09246_ (.A1(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_en ),
    .A2(clknet_3_6__leaf__00564_),
    .ZN(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ));
 AND2_X1 _09247_ (.A1(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_en ),
    .A2(clknet_3_6__leaf__00564_),
    .ZN(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ));
 AND2_X1 _09248_ (.A1(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_en ),
    .A2(clknet_3_4__leaf__00564_),
    .ZN(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ));
 AND2_X1 _09249_ (.A1(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_en ),
    .A2(clknet_3_2__leaf__00564_),
    .ZN(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ));
 AND2_X1 _09250_ (.A1(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_en ),
    .A2(clknet_3_6__leaf__00564_),
    .ZN(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ));
 AND2_X1 _09251_ (.A1(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_en ),
    .A2(clknet_3_2__leaf__00564_),
    .ZN(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ));
 AND2_X1 _09252_ (.A1(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_en ),
    .A2(clknet_3_5__leaf__00564_),
    .ZN(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ));
 AND2_X1 _09253_ (.A1(\lut.gen_sub_units_scm.__4.sub_unit_i.cg_we_global.clk_en ),
    .A2(clknet_2_1__leaf__00532_),
    .ZN(_00567_));
 TAPCELL_X1 PHY_21 ();
 AND2_X1 _09255_ (.A1(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_en ),
    .A2(clknet_3_4__leaf__00567_),
    .ZN(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ));
 AND2_X1 _09256_ (.A1(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_en ),
    .A2(clknet_3_1__leaf__00567_),
    .ZN(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ));
 AND2_X1 _09257_ (.A1(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_en ),
    .A2(clknet_3_0__leaf__00567_),
    .ZN(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ));
 AND2_X1 _09258_ (.A1(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_en ),
    .A2(clknet_3_7__leaf__00567_),
    .ZN(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ));
 AND2_X1 _09259_ (.A1(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_en ),
    .A2(clknet_3_2__leaf__00567_),
    .ZN(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ));
 AND2_X1 _09260_ (.A1(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_en ),
    .A2(clknet_3_0__leaf__00567_),
    .ZN(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ));
 AND2_X1 _09261_ (.A1(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_en ),
    .A2(clknet_3_7__leaf__00567_),
    .ZN(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ));
 AND2_X1 _09262_ (.A1(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_en ),
    .A2(clknet_3_5__leaf__00567_),
    .ZN(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ));
 AND2_X1 _09263_ (.A1(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_en ),
    .A2(clknet_3_2__leaf__00567_),
    .ZN(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ));
 TAPCELL_X1 PHY_20 ();
 AND2_X1 _09265_ (.A1(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_en ),
    .A2(clknet_3_2__leaf__00567_),
    .ZN(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ));
 AND2_X1 _09266_ (.A1(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_en ),
    .A2(clknet_3_1__leaf__00567_),
    .ZN(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ));
 AND2_X1 _09267_ (.A1(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_en ),
    .A2(clknet_3_2__leaf__00567_),
    .ZN(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ));
 AND2_X1 _09268_ (.A1(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_en ),
    .A2(clknet_3_0__leaf__00567_),
    .ZN(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ));
 AND2_X1 _09269_ (.A1(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_en ),
    .A2(clknet_3_6__leaf__00567_),
    .ZN(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ));
 AND2_X1 _09270_ (.A1(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_en ),
    .A2(clknet_3_1__leaf__00567_),
    .ZN(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ));
 AND2_X1 _09271_ (.A1(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_en ),
    .A2(clknet_3_6__leaf__00567_),
    .ZN(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ));
 AND2_X1 _09272_ (.A1(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_en ),
    .A2(clknet_3_5__leaf__00567_),
    .ZN(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ));
 AND2_X1 _09273_ (.A1(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_en ),
    .A2(clknet_3_7__leaf__00567_),
    .ZN(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ));
 AND2_X1 _09274_ (.A1(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_en ),
    .A2(clknet_3_6__leaf__00567_),
    .ZN(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ));
 TAPCELL_X1 PHY_19 ();
 AND2_X1 _09276_ (.A1(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_en ),
    .A2(clknet_3_5__leaf__00567_),
    .ZN(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ));
 AND2_X1 _09277_ (.A1(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_en ),
    .A2(clknet_3_7__leaf__00567_),
    .ZN(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ));
 AND2_X1 _09278_ (.A1(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_en ),
    .A2(clknet_3_3__leaf__00567_),
    .ZN(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ));
 AND2_X1 _09279_ (.A1(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_en ),
    .A2(clknet_3_5__leaf__00567_),
    .ZN(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ));
 AND2_X1 _09280_ (.A1(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_en ),
    .A2(clknet_3_7__leaf__00567_),
    .ZN(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ));
 AND2_X1 _09281_ (.A1(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_en ),
    .A2(clknet_3_1__leaf__00567_),
    .ZN(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ));
 AND2_X1 _09282_ (.A1(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_en ),
    .A2(clknet_3_3__leaf__00567_),
    .ZN(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ));
 AND2_X1 _09283_ (.A1(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_en ),
    .A2(clknet_3_0__leaf__00567_),
    .ZN(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ));
 AND2_X1 _09284_ (.A1(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_en ),
    .A2(clknet_3_1__leaf__00567_),
    .ZN(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ));
 AND2_X1 _09285_ (.A1(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_en ),
    .A2(clknet_3_7__leaf__00567_),
    .ZN(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ));
 AND2_X1 _09286_ (.A1(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_en ),
    .A2(clknet_3_4__leaf__00567_),
    .ZN(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ));
 AND2_X1 _09287_ (.A1(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_en ),
    .A2(clknet_3_4__leaf__00567_),
    .ZN(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ));
 AND2_X1 _09288_ (.A1(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_en ),
    .A2(clknet_3_2__leaf__00567_),
    .ZN(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ));
 AND2_X1 _09289_ (.A1(\lut.gen_sub_units_scm.__3.sub_unit_i.cg_we_global.clk_en ),
    .A2(clknet_2_2__leaf__00532_),
    .ZN(_00570_));
 TAPCELL_X1 PHY_18 ();
 AND2_X1 _09291_ (.A1(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_en ),
    .A2(clknet_3_7__leaf__00570_),
    .ZN(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ));
 AND2_X1 _09292_ (.A1(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_en ),
    .A2(clknet_3_0__leaf__00570_),
    .ZN(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ));
 AND2_X1 _09293_ (.A1(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_en ),
    .A2(clknet_3_3__leaf__00570_),
    .ZN(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ));
 AND2_X1 _09294_ (.A1(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_en ),
    .A2(clknet_3_1__leaf__00570_),
    .ZN(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ));
 AND2_X1 _09295_ (.A1(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_en ),
    .A2(clknet_3_2__leaf__00570_),
    .ZN(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ));
 AND2_X1 _09296_ (.A1(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_en ),
    .A2(clknet_3_5__leaf__00570_),
    .ZN(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ));
 AND2_X1 _09297_ (.A1(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_en ),
    .A2(clknet_3_6__leaf__00570_),
    .ZN(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ));
 AND2_X1 _09298_ (.A1(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_en ),
    .A2(clknet_3_7__leaf__00570_),
    .ZN(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ));
 AND2_X1 _09299_ (.A1(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_en ),
    .A2(clknet_3_6__leaf__00570_),
    .ZN(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ));
 TAPCELL_X1 PHY_17 ();
 AND2_X1 _09301_ (.A1(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_en ),
    .A2(clknet_3_6__leaf__00570_),
    .ZN(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ));
 AND2_X1 _09302_ (.A1(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_en ),
    .A2(clknet_3_7__leaf__00570_),
    .ZN(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ));
 AND2_X1 _09303_ (.A1(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_en ),
    .A2(clknet_3_6__leaf__00570_),
    .ZN(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ));
 AND2_X1 _09304_ (.A1(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_en ),
    .A2(clknet_3_3__leaf__00570_),
    .ZN(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ));
 AND2_X1 _09305_ (.A1(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_en ),
    .A2(clknet_3_0__leaf__00570_),
    .ZN(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ));
 AND2_X1 _09306_ (.A1(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_en ),
    .A2(clknet_3_1__leaf__00570_),
    .ZN(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ));
 AND2_X1 _09307_ (.A1(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_en ),
    .A2(clknet_3_2__leaf__00570_),
    .ZN(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ));
 AND2_X1 _09308_ (.A1(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_en ),
    .A2(clknet_3_1__leaf__00570_),
    .ZN(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ));
 AND2_X1 _09309_ (.A1(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_en ),
    .A2(clknet_3_1__leaf__00570_),
    .ZN(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ));
 AND2_X1 _09310_ (.A1(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_en ),
    .A2(clknet_3_2__leaf__00570_),
    .ZN(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ));
 TAPCELL_X1 PHY_16 ();
 AND2_X1 _09312_ (.A1(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_en ),
    .A2(clknet_3_2__leaf__00570_),
    .ZN(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ));
 AND2_X1 _09313_ (.A1(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_en ),
    .A2(clknet_3_4__leaf__00570_),
    .ZN(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ));
 AND2_X1 _09314_ (.A1(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_en ),
    .A2(clknet_3_4__leaf__00570_),
    .ZN(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ));
 AND2_X1 _09315_ (.A1(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_en ),
    .A2(clknet_3_0__leaf__00570_),
    .ZN(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ));
 AND2_X1 _09316_ (.A1(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_en ),
    .A2(clknet_3_4__leaf__00570_),
    .ZN(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ));
 AND2_X1 _09317_ (.A1(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_en ),
    .A2(clknet_3_5__leaf__00570_),
    .ZN(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ));
 AND2_X1 _09318_ (.A1(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_en ),
    .A2(clknet_3_6__leaf__00570_),
    .ZN(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ));
 AND2_X1 _09319_ (.A1(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_en ),
    .A2(clknet_3_1__leaf__00570_),
    .ZN(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ));
 AND2_X1 _09320_ (.A1(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_en ),
    .A2(clknet_3_5__leaf__00570_),
    .ZN(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ));
 AND2_X1 _09321_ (.A1(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_en ),
    .A2(clknet_3_5__leaf__00570_),
    .ZN(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ));
 AND2_X1 _09322_ (.A1(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_en ),
    .A2(clknet_3_5__leaf__00570_),
    .ZN(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ));
 AND2_X1 _09323_ (.A1(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_en ),
    .A2(clknet_3_3__leaf__00570_),
    .ZN(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ));
 AND2_X1 _09324_ (.A1(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_en ),
    .A2(clknet_3_7__leaf__00570_),
    .ZN(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ));
 AND2_X1 _09325_ (.A1(\lut.gen_sub_units_scm.__2.sub_unit_i.cg_we_global.clk_en ),
    .A2(clknet_2_2__leaf__00532_),
    .ZN(_00573_));
 TAPCELL_X1 PHY_15 ();
 AND2_X1 _09327_ (.A1(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_en ),
    .A2(clknet_3_2__leaf__00573_),
    .ZN(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ));
 AND2_X1 _09328_ (.A1(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_en ),
    .A2(clknet_3_5__leaf__00573_),
    .ZN(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ));
 AND2_X1 _09329_ (.A1(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_en ),
    .A2(clknet_3_5__leaf__00573_),
    .ZN(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ));
 AND2_X1 _09330_ (.A1(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_en ),
    .A2(clknet_3_0__leaf__00573_),
    .ZN(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ));
 AND2_X1 _09331_ (.A1(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_en ),
    .A2(clknet_3_7__leaf__00573_),
    .ZN(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ));
 AND2_X1 _09332_ (.A1(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_en ),
    .A2(clknet_3_6__leaf__00573_),
    .ZN(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ));
 AND2_X1 _09333_ (.A1(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_en ),
    .A2(clknet_3_6__leaf__00573_),
    .ZN(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ));
 AND2_X1 _09334_ (.A1(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_en ),
    .A2(clknet_3_1__leaf__00573_),
    .ZN(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ));
 AND2_X1 _09335_ (.A1(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_en ),
    .A2(clknet_3_0__leaf__00573_),
    .ZN(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ));
 TAPCELL_X1 PHY_14 ();
 AND2_X1 _09337_ (.A1(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_en ),
    .A2(clknet_3_7__leaf__00573_),
    .ZN(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ));
 AND2_X1 _09338_ (.A1(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_en ),
    .A2(clknet_3_7__leaf__00573_),
    .ZN(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ));
 AND2_X1 _09339_ (.A1(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_en ),
    .A2(clknet_3_7__leaf__00573_),
    .ZN(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ));
 AND2_X1 _09340_ (.A1(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_en ),
    .A2(clknet_3_5__leaf__00573_),
    .ZN(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ));
 AND2_X1 _09341_ (.A1(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_en ),
    .A2(clknet_3_5__leaf__00573_),
    .ZN(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ));
 AND2_X1 _09342_ (.A1(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_en ),
    .A2(clknet_3_5__leaf__00573_),
    .ZN(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ));
 AND2_X1 _09343_ (.A1(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_en ),
    .A2(clknet_3_1__leaf__00573_),
    .ZN(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ));
 AND2_X1 _09344_ (.A1(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_en ),
    .A2(clknet_3_1__leaf__00573_),
    .ZN(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ));
 AND2_X1 _09345_ (.A1(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_en ),
    .A2(clknet_3_3__leaf__00573_),
    .ZN(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ));
 AND2_X1 _09346_ (.A1(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_en ),
    .A2(clknet_3_5__leaf__00573_),
    .ZN(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ));
 TAPCELL_X1 PHY_13 ();
 AND2_X1 _09348_ (.A1(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_en ),
    .A2(clknet_3_4__leaf__00573_),
    .ZN(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ));
 AND2_X1 _09349_ (.A1(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_en ),
    .A2(clknet_3_7__leaf__00573_),
    .ZN(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ));
 AND2_X1 _09350_ (.A1(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_en ),
    .A2(clknet_3_2__leaf__00573_),
    .ZN(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ));
 AND2_X1 _09351_ (.A1(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_en ),
    .A2(clknet_3_4__leaf__00573_),
    .ZN(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ));
 AND2_X1 _09352_ (.A1(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_en ),
    .A2(clknet_3_3__leaf__00573_),
    .ZN(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ));
 AND2_X1 _09353_ (.A1(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_en ),
    .A2(clknet_3_3__leaf__00573_),
    .ZN(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ));
 AND2_X1 _09354_ (.A1(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_en ),
    .A2(clknet_3_6__leaf__00573_),
    .ZN(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ));
 AND2_X1 _09355_ (.A1(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_en ),
    .A2(clknet_3_3__leaf__00573_),
    .ZN(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ));
 AND2_X1 _09356_ (.A1(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_en ),
    .A2(clknet_3_3__leaf__00573_),
    .ZN(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ));
 AND2_X1 _09357_ (.A1(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_en ),
    .A2(clknet_3_2__leaf__00573_),
    .ZN(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ));
 AND2_X1 _09358_ (.A1(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_en ),
    .A2(clknet_3_3__leaf__00573_),
    .ZN(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ));
 AND2_X1 _09359_ (.A1(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_en ),
    .A2(clknet_3_6__leaf__00573_),
    .ZN(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ));
 AND2_X1 _09360_ (.A1(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_en ),
    .A2(clknet_3_7__leaf__00573_),
    .ZN(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ));
 AND2_X1 _09361_ (.A1(\lut.gen_sub_units_scm.__1.sub_unit_i.cg_we_global.clk_en ),
    .A2(clknet_2_3__leaf__00532_),
    .ZN(_00576_));
 TAPCELL_X1 PHY_12 ();
 AND2_X1 _09363_ (.A1(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_en ),
    .A2(clknet_3_1__leaf__00576_),
    .ZN(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ));
 AND2_X1 _09364_ (.A1(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_en ),
    .A2(clknet_3_6__leaf__00576_),
    .ZN(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ));
 AND2_X1 _09365_ (.A1(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_en ),
    .A2(clknet_3_0__leaf__00576_),
    .ZN(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ));
 AND2_X1 _09366_ (.A1(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_en ),
    .A2(clknet_3_6__leaf__00576_),
    .ZN(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ));
 AND2_X1 _09367_ (.A1(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_en ),
    .A2(clknet_3_7__leaf__00576_),
    .ZN(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ));
 AND2_X1 _09368_ (.A1(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_en ),
    .A2(clknet_3_6__leaf__00576_),
    .ZN(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ));
 AND2_X1 _09369_ (.A1(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_en ),
    .A2(clknet_3_7__leaf__00576_),
    .ZN(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ));
 AND2_X1 _09370_ (.A1(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_en ),
    .A2(clknet_3_5__leaf__00576_),
    .ZN(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ));
 AND2_X1 _09371_ (.A1(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_en ),
    .A2(clknet_3_5__leaf__00576_),
    .ZN(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ));
 TAPCELL_X1 PHY_11 ();
 AND2_X1 _09373_ (.A1(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_en ),
    .A2(clknet_3_2__leaf__00576_),
    .ZN(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ));
 AND2_X1 _09374_ (.A1(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_en ),
    .A2(clknet_3_2__leaf__00576_),
    .ZN(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ));
 AND2_X1 _09375_ (.A1(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_en ),
    .A2(clknet_3_7__leaf__00576_),
    .ZN(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ));
 AND2_X1 _09376_ (.A1(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_en ),
    .A2(clknet_3_1__leaf__00576_),
    .ZN(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ));
 AND2_X1 _09377_ (.A1(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_en ),
    .A2(clknet_3_4__leaf__00576_),
    .ZN(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ));
 AND2_X1 _09378_ (.A1(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_en ),
    .A2(clknet_3_1__leaf__00576_),
    .ZN(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ));
 AND2_X1 _09379_ (.A1(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_en ),
    .A2(clknet_3_4__leaf__00576_),
    .ZN(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ));
 AND2_X1 _09380_ (.A1(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_en ),
    .A2(clknet_3_3__leaf__00576_),
    .ZN(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ));
 AND2_X1 _09381_ (.A1(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_en ),
    .A2(clknet_3_6__leaf__00576_),
    .ZN(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ));
 AND2_X1 _09382_ (.A1(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_en ),
    .A2(clknet_3_2__leaf__00576_),
    .ZN(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ));
 TAPCELL_X1 PHY_10 ();
 AND2_X1 _09384_ (.A1(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_en ),
    .A2(clknet_3_3__leaf__00576_),
    .ZN(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ));
 AND2_X1 _09385_ (.A1(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_en ),
    .A2(clknet_3_4__leaf__00576_),
    .ZN(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ));
 AND2_X1 _09386_ (.A1(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_en ),
    .A2(clknet_3_6__leaf__00576_),
    .ZN(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ));
 AND2_X1 _09387_ (.A1(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_en ),
    .A2(clknet_3_2__leaf__00576_),
    .ZN(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ));
 AND2_X1 _09388_ (.A1(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_en ),
    .A2(clknet_3_3__leaf__00576_),
    .ZN(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ));
 AND2_X1 _09389_ (.A1(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_en ),
    .A2(clknet_3_5__leaf__00576_),
    .ZN(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ));
 AND2_X1 _09390_ (.A1(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_en ),
    .A2(clknet_3_3__leaf__00576_),
    .ZN(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ));
 AND2_X1 _09391_ (.A1(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_en ),
    .A2(clknet_3_0__leaf__00576_),
    .ZN(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ));
 AND2_X1 _09392_ (.A1(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_en ),
    .A2(clknet_3_7__leaf__00576_),
    .ZN(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ));
 AND2_X1 _09393_ (.A1(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_en ),
    .A2(clknet_3_7__leaf__00576_),
    .ZN(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ));
 AND2_X1 _09394_ (.A1(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_en ),
    .A2(clknet_3_7__leaf__00576_),
    .ZN(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ));
 AND2_X1 _09395_ (.A1(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_en ),
    .A2(clknet_3_7__leaf__00576_),
    .ZN(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ));
 AND2_X1 _09396_ (.A1(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_en ),
    .A2(clknet_3_4__leaf__00576_),
    .ZN(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ));
 AND2_X1 _09397_ (.A1(\lut.gen_sub_units_scm.__0.sub_unit_i.cg_we_global.clk_en ),
    .A2(clknet_2_3__leaf__00532_),
    .ZN(_00579_));
 TAPCELL_X1 PHY_9 ();
 AND2_X1 _09399_ (.A1(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_en ),
    .A2(clknet_3_4__leaf__00579_),
    .ZN(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ));
 AND2_X1 _09400_ (.A1(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_en ),
    .A2(clknet_3_0__leaf__00579_),
    .ZN(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ));
 AND2_X1 _09401_ (.A1(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_en ),
    .A2(clknet_3_1__leaf__00579_),
    .ZN(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ));
 AND2_X1 _09402_ (.A1(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_en ),
    .A2(clknet_3_6__leaf__00579_),
    .ZN(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ));
 AND2_X1 _09403_ (.A1(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_en ),
    .A2(clknet_3_2__leaf__00579_),
    .ZN(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ));
 AND2_X1 _09404_ (.A1(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_en ),
    .A2(clknet_3_0__leaf__00579_),
    .ZN(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ));
 AND2_X1 _09405_ (.A1(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_en ),
    .A2(clknet_3_4__leaf__00579_),
    .ZN(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ));
 AND2_X1 _09406_ (.A1(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_en ),
    .A2(clknet_3_7__leaf__00579_),
    .ZN(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ));
 AND2_X1 _09407_ (.A1(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_en ),
    .A2(clknet_3_6__leaf__00579_),
    .ZN(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ));
 TAPCELL_X1 PHY_8 ();
 AND2_X1 _09409_ (.A1(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_en ),
    .A2(clknet_3_7__leaf__00579_),
    .ZN(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ));
 AND2_X1 _09410_ (.A1(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_en ),
    .A2(clknet_3_6__leaf__00579_),
    .ZN(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ));
 AND2_X1 _09411_ (.A1(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_en ),
    .A2(clknet_3_2__leaf__00579_),
    .ZN(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ));
 AND2_X1 _09412_ (.A1(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_en ),
    .A2(clknet_3_1__leaf__00579_),
    .ZN(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ));
 AND2_X1 _09413_ (.A1(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_en ),
    .A2(clknet_3_6__leaf__00579_),
    .ZN(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ));
 AND2_X1 _09414_ (.A1(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_en ),
    .A2(clknet_3_7__leaf__00579_),
    .ZN(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ));
 AND2_X1 _09415_ (.A1(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_en ),
    .A2(clknet_3_2__leaf__00579_),
    .ZN(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ));
 AND2_X1 _09416_ (.A1(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_en ),
    .A2(clknet_3_5__leaf__00579_),
    .ZN(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ));
 AND2_X1 _09417_ (.A1(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_en ),
    .A2(clknet_3_7__leaf__00579_),
    .ZN(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ));
 AND2_X1 _09418_ (.A1(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_en ),
    .A2(clknet_3_5__leaf__00579_),
    .ZN(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ));
 TAPCELL_X1 PHY_7 ();
 AND2_X1 _09420_ (.A1(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_en ),
    .A2(clknet_3_5__leaf__00579_),
    .ZN(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ));
 AND2_X1 _09421_ (.A1(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_en ),
    .A2(clknet_3_7__leaf__00579_),
    .ZN(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ));
 AND2_X1 _09422_ (.A1(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_en ),
    .A2(clknet_3_3__leaf__00579_),
    .ZN(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ));
 AND2_X1 _09423_ (.A1(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_en ),
    .A2(clknet_3_1__leaf__00579_),
    .ZN(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ));
 AND2_X1 _09424_ (.A1(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_en ),
    .A2(clknet_3_2__leaf__00579_),
    .ZN(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ));
 AND2_X1 _09425_ (.A1(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_en ),
    .A2(clknet_3_4__leaf__00579_),
    .ZN(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ));
 AND2_X1 _09426_ (.A1(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_en ),
    .A2(clknet_3_6__leaf__00579_),
    .ZN(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ));
 AND2_X1 _09427_ (.A1(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_en ),
    .A2(clknet_3_6__leaf__00579_),
    .ZN(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ));
 AND2_X1 _09428_ (.A1(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_en ),
    .A2(clknet_3_6__leaf__00579_),
    .ZN(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ));
 AND2_X1 _09429_ (.A1(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_en ),
    .A2(clknet_3_1__leaf__00579_),
    .ZN(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ));
 AND2_X1 _09430_ (.A1(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_en ),
    .A2(clknet_3_1__leaf__00579_),
    .ZN(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ));
 AND2_X1 _09431_ (.A1(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_en ),
    .A2(clknet_3_3__leaf__00579_),
    .ZN(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ));
 AND2_X1 _09432_ (.A1(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_en ),
    .A2(clknet_3_5__leaf__00579_),
    .ZN(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ));
 NOR2_X1 _09433_ (.A1(_00870_),
    .A2(_00897_),
    .ZN(_00582_));
 NOR2_X1 _09434_ (.A1(_00582_),
    .A2(_00895_),
    .ZN(_04239_));
 INV_X1 _09435_ (.A(_00903_),
    .ZN(_04243_));
 NAND2_X1 _09436_ (.A1(_04293_),
    .A2(_04291_),
    .ZN(_00583_));
 OAI21_X1 _09437_ (.A(_00890_),
    .B1(_00583_),
    .B2(_04232_),
    .ZN(_04236_));
 MUX2_X1 _09438_ (.A(_04253_),
    .B(net30),
    .S(_00827_),
    .Z(_00584_));
 AND2_X1 _09439_ (.A1(net6),
    .A2(_00584_),
    .ZN(_00000_));
 TAPCELL_X1 PHY_6 ();
 NOR2_X1 _09441_ (.A1(_04198_),
    .A2(_00827_),
    .ZN(_00586_));
 TAPCELL_X1 PHY_5 ();
 AOI21_X1 _09443_ (.A(_00586_),
    .B1(_00827_),
    .B2(net41),
    .ZN(_00588_));
 NOR2_X1 _09444_ (.A1(_00907_),
    .A2(_00588_),
    .ZN(_00001_));
 MUX2_X1 _09445_ (.A(_04200_),
    .B(net52),
    .S(_00827_),
    .Z(_00589_));
 AND2_X1 _09446_ (.A1(net6),
    .A2(_00589_),
    .ZN(_00002_));
 TAPCELL_X1 PHY_4 ();
 TAPCELL_X1 PHY_3 ();
 OR2_X1 _09449_ (.A1(_00827_),
    .A2(_00834_),
    .ZN(_00592_));
 TAPCELL_X1 PHY_2 ();
 NAND2_X1 _09451_ (.A1(net55),
    .A2(_00827_),
    .ZN(_00594_));
 AOI21_X1 _09452_ (.A(_00907_),
    .B1(_00592_),
    .B2(_00594_),
    .ZN(_00003_));
 MUX2_X1 _09453_ (.A(_04203_),
    .B(net56),
    .S(_00827_),
    .Z(_00595_));
 AND2_X1 _09454_ (.A1(net6),
    .A2(_00595_),
    .ZN(_00004_));
 OR2_X1 _09455_ (.A1(_00827_),
    .A2(_00838_),
    .ZN(_00596_));
 NAND2_X1 _09456_ (.A1(net57),
    .A2(_00827_),
    .ZN(_00597_));
 AOI21_X1 _09457_ (.A(_00907_),
    .B1(_00596_),
    .B2(_00597_),
    .ZN(_00005_));
 NOR2_X1 _09458_ (.A1(_04208_),
    .A2(_00827_),
    .ZN(_00598_));
 AOI21_X1 _09459_ (.A(_00598_),
    .B1(_00827_),
    .B2(net58),
    .ZN(_00599_));
 NOR2_X1 _09460_ (.A1(_00907_),
    .A2(_00599_),
    .ZN(_00006_));
 OR2_X1 _09461_ (.A1(_00827_),
    .A2(_00844_),
    .ZN(_00600_));
 NAND2_X1 _09462_ (.A1(net59),
    .A2(_00827_),
    .ZN(_00601_));
 AOI21_X1 _09463_ (.A(_00907_),
    .B1(_00600_),
    .B2(_00601_),
    .ZN(_00007_));
 MUX2_X1 _09464_ (.A(_04211_),
    .B(net60),
    .S(_00827_),
    .Z(_00602_));
 AND2_X1 _09465_ (.A1(net6),
    .A2(_00602_),
    .ZN(_00008_));
 TAPCELL_X1 PHY_1 ();
 TAPCELL_X1 PHY_0 ();
 OR2_X1 _09468_ (.A1(_00827_),
    .A2(_00848_),
    .ZN(_00605_));
 NAND2_X1 _09469_ (.A1(net61),
    .A2(_00827_),
    .ZN(_00606_));
 AOI21_X1 _09470_ (.A(_00907_),
    .B1(_00605_),
    .B2(_00606_),
    .ZN(_00009_));
 NOR2_X1 _09471_ (.A1(_04216_),
    .A2(_00827_),
    .ZN(_00607_));
 AOI21_X1 _09472_ (.A(_00607_),
    .B1(_00827_),
    .B2(net31),
    .ZN(_00608_));
 NOR2_X1 _09473_ (.A1(_00907_),
    .A2(_00608_),
    .ZN(_00010_));
 OR2_X1 _09474_ (.A1(_00827_),
    .A2(_00852_),
    .ZN(_00609_));
 NAND2_X1 _09475_ (.A1(net32),
    .A2(_00827_),
    .ZN(_00610_));
 AOI21_X1 _09476_ (.A(_00907_),
    .B1(_00609_),
    .B2(_00610_),
    .ZN(_00011_));
 NOR2_X1 _09477_ (.A1(_04220_),
    .A2(_00827_),
    .ZN(_00611_));
 AOI21_X1 _09478_ (.A(_00611_),
    .B1(_00827_),
    .B2(net33),
    .ZN(_00612_));
 NOR2_X1 _09479_ (.A1(_00907_),
    .A2(_00612_),
    .ZN(_00012_));
 OR2_X1 _09480_ (.A1(_00827_),
    .A2(_00862_),
    .ZN(_00613_));
 NAND2_X1 _09481_ (.A1(net34),
    .A2(_00827_),
    .ZN(_00614_));
 AOI21_X1 _09482_ (.A(_00907_),
    .B1(_00613_),
    .B2(_00614_),
    .ZN(_00013_));
 NOR2_X1 _09483_ (.A1(_04224_),
    .A2(_00827_),
    .ZN(_00615_));
 AOI21_X1 _09484_ (.A(_00615_),
    .B1(_00827_),
    .B2(net35),
    .ZN(_00616_));
 NOR2_X1 _09485_ (.A1(_00907_),
    .A2(_00616_),
    .ZN(_00014_));
 OR2_X1 _09486_ (.A1(_00827_),
    .A2(_00865_),
    .ZN(_00617_));
 NAND2_X1 _09487_ (.A1(net36),
    .A2(_00827_),
    .ZN(_00618_));
 AOI21_X1 _09488_ (.A(_00907_),
    .B1(_00617_),
    .B2(_00618_),
    .ZN(_00015_));
 MUX2_X1 _09489_ (.A(_04227_),
    .B(net37),
    .S(_00827_),
    .Z(_00619_));
 AND2_X1 _09490_ (.A1(net6),
    .A2(_00619_),
    .ZN(_00016_));
 OR2_X1 _09491_ (.A1(_00827_),
    .A2(_00871_),
    .ZN(_00620_));
 NAND2_X1 _09492_ (.A1(net38),
    .A2(_00827_),
    .ZN(_00621_));
 AOI21_X1 _09493_ (.A(_00907_),
    .B1(_00620_),
    .B2(_00621_),
    .ZN(_00017_));
 NOR2_X1 _09494_ (.A1(_04231_),
    .A2(_00827_),
    .ZN(_00622_));
 AOI21_X1 _09495_ (.A(_00622_),
    .B1(_00827_),
    .B2(net39),
    .ZN(_00623_));
 NOR2_X1 _09496_ (.A1(_00907_),
    .A2(_00623_),
    .ZN(_00018_));
 OR2_X1 _09497_ (.A1(_00827_),
    .A2(_00873_),
    .ZN(_00624_));
 NAND2_X1 _09498_ (.A1(net40),
    .A2(_00827_),
    .ZN(_00625_));
 AOI21_X1 _09499_ (.A(_00907_),
    .B1(_00624_),
    .B2(_00625_),
    .ZN(_00019_));
 NOR2_X1 _09500_ (.A1(_04235_),
    .A2(_00827_),
    .ZN(_00626_));
 AOI21_X1 _09501_ (.A(_00626_),
    .B1(_00827_),
    .B2(net42),
    .ZN(_00627_));
 NOR2_X1 _09502_ (.A1(_00907_),
    .A2(_00627_),
    .ZN(_00020_));
 OR2_X1 _09503_ (.A1(_00827_),
    .A2(_00882_),
    .ZN(_00628_));
 NAND2_X1 _09504_ (.A1(net43),
    .A2(_00827_),
    .ZN(_00629_));
 AOI21_X1 _09505_ (.A(_00907_),
    .B1(_00628_),
    .B2(_00629_),
    .ZN(_00021_));
 NOR2_X1 _09506_ (.A1(_04238_),
    .A2(_00827_),
    .ZN(_00630_));
 AOI21_X1 _09507_ (.A(_00630_),
    .B1(_00827_),
    .B2(net44),
    .ZN(_00631_));
 NOR2_X1 _09508_ (.A1(_00907_),
    .A2(_00631_),
    .ZN(_00022_));
 OR2_X1 _09509_ (.A1(_00827_),
    .A2(_00883_),
    .ZN(_00632_));
 NAND2_X1 _09510_ (.A1(net45),
    .A2(_00827_),
    .ZN(_00633_));
 AOI21_X1 _09511_ (.A(_00907_),
    .B1(_00632_),
    .B2(_00633_),
    .ZN(_00023_));
 MUX2_X1 _09512_ (.A(_04242_),
    .B(net46),
    .S(_00827_),
    .Z(_00634_));
 AND2_X1 _09513_ (.A1(net6),
    .A2(_00634_),
    .ZN(_00024_));
 OR2_X1 _09514_ (.A1(_00827_),
    .A2(_00884_),
    .ZN(_00635_));
 NAND2_X1 _09515_ (.A1(net47),
    .A2(_00827_),
    .ZN(_00636_));
 AOI21_X1 _09516_ (.A(_00907_),
    .B1(_00635_),
    .B2(_00636_),
    .ZN(_00025_));
 NOR2_X1 _09517_ (.A1(_04245_),
    .A2(_00827_),
    .ZN(_00637_));
 AOI21_X1 _09518_ (.A(_00637_),
    .B1(_00827_),
    .B2(net48),
    .ZN(_00638_));
 NOR2_X1 _09519_ (.A1(_00907_),
    .A2(_00638_),
    .ZN(_00026_));
 OR2_X1 _09520_ (.A1(_00827_),
    .A2(_00885_),
    .ZN(_00639_));
 NAND2_X1 _09521_ (.A1(net49),
    .A2(_00827_),
    .ZN(_00640_));
 AOI21_X1 _09522_ (.A(_00907_),
    .B1(_00639_),
    .B2(_00640_),
    .ZN(_00027_));
 NOR2_X1 _09523_ (.A1(_04248_),
    .A2(_00827_),
    .ZN(_00641_));
 AOI21_X1 _09524_ (.A(_00641_),
    .B1(_00827_),
    .B2(net50),
    .ZN(_00642_));
 NOR2_X1 _09525_ (.A1(_00907_),
    .A2(_00642_),
    .ZN(_00028_));
 OR2_X1 _09526_ (.A1(_00827_),
    .A2(_00886_),
    .ZN(_00643_));
 NAND2_X1 _09527_ (.A1(net51),
    .A2(_00827_),
    .ZN(_00644_));
 AOI21_X1 _09528_ (.A(_00907_),
    .B1(_00643_),
    .B2(_00644_),
    .ZN(_00029_));
 NOR2_X1 _09529_ (.A1(_04252_),
    .A2(_00827_),
    .ZN(_00645_));
 AOI21_X1 _09530_ (.A(_00645_),
    .B1(_00827_),
    .B2(net53),
    .ZN(_00646_));
 NOR2_X1 _09531_ (.A1(_00907_),
    .A2(_00646_),
    .ZN(_00030_));
 NOR2_X1 _09532_ (.A1(_00827_),
    .A2(_00906_),
    .ZN(_00647_));
 AOI21_X1 _09533_ (.A(_00647_),
    .B1(_00827_),
    .B2(net54),
    .ZN(_00648_));
 NOR2_X1 _09534_ (.A1(_00907_),
    .A2(_00648_),
    .ZN(_00031_));
 MUX2_X1 _09535_ (.A(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[0] ),
    .B(net21),
    .S(net29),
    .Z(_00032_));
 MUX2_X1 _09536_ (.A(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[1] ),
    .B(net22),
    .S(net29),
    .Z(_00033_));
 MUX2_X1 _09537_ (.A(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[2] ),
    .B(net23),
    .S(net29),
    .Z(_00034_));
 MUX2_X1 _09538_ (.A(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[3] ),
    .B(net24),
    .S(net29),
    .Z(_00035_));
 MUX2_X1 _09539_ (.A(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[4] ),
    .B(net25),
    .S(net29),
    .Z(_00036_));
 MUX2_X1 _09540_ (.A(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[5] ),
    .B(net26),
    .S(net29),
    .Z(_00037_));
 MUX2_X1 _09541_ (.A(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[6] ),
    .B(net27),
    .S(net29),
    .Z(_00038_));
 MUX2_X1 _09542_ (.A(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[7] ),
    .B(net28),
    .S(net29),
    .Z(_00039_));
 NOR4_X1 _09543_ (.A1(\caddr_q[1] ),
    .A2(\caddr_q[0] ),
    .A3(\caddr_q[3] ),
    .A4(\caddr_q[2] ),
    .ZN(_00649_));
 NAND3_X1 _09544_ (.A1(_00825_),
    .A2(net62),
    .A3(_00649_),
    .ZN(_00650_));
 AOI21_X1 _09545_ (.A(_00907_),
    .B1(_00827_),
    .B2(_00650_),
    .ZN(_00040_));
 FA_X1 _09546_ (.A(_04196_),
    .B(\genblk1.gen_int_accumulation.int_adder.int_short_converted[1] ),
    .CI(\genblk1.gen_int_accumulation.int_adder.int_long_i[1] ),
    .CO(_04197_),
    .S(_04198_));
 FA_X1 _09547_ (.A(_04197_),
    .B(\genblk1.gen_int_accumulation.int_adder.int_short_converted[2] ),
    .CI(\genblk1.gen_int_accumulation.int_adder.int_long_i[2] ),
    .CO(_04199_),
    .S(_04200_));
 FA_X1 _09548_ (.A(_04201_),
    .B(\genblk1.gen_int_accumulation.int_adder.int_short_converted[4] ),
    .CI(\genblk1.gen_int_accumulation.int_adder.int_long_i[4] ),
    .CO(_04202_),
    .S(_04203_));
 FA_X1 _09549_ (.A(_04204_),
    .B(_04205_),
    .CI(_04206_),
    .CO(_04207_),
    .S(_04208_));
 FA_X1 _09550_ (.A(_04209_),
    .B(\genblk1.gen_int_accumulation.int_adder.int_short_converted[10] ),
    .CI(\genblk1.gen_int_accumulation.int_adder.int_long_i[8] ),
    .CO(_04210_),
    .S(_04211_));
 FA_X1 _09551_ (.A(_04212_),
    .B(_04213_),
    .CI(_04214_),
    .CO(_04215_),
    .S(_04216_));
 FA_X1 _09552_ (.A(_04217_),
    .B(_04213_),
    .CI(_04218_),
    .CO(_04219_),
    .S(_04220_));
 FA_X1 _09553_ (.A(_04221_),
    .B(_04213_),
    .CI(_04222_),
    .CO(_04223_),
    .S(_04224_));
 FA_X1 _09554_ (.A(_04225_),
    .B(\genblk1.gen_int_accumulation.int_adder.int_short_converted[10] ),
    .CI(\genblk1.gen_int_accumulation.int_adder.int_long_i[16] ),
    .CO(_04226_),
    .S(_04227_));
 FA_X1 _09555_ (.A(_04228_),
    .B(_04213_),
    .CI(_04229_),
    .CO(_04230_),
    .S(_04231_));
 FA_X1 _09556_ (.A(_04232_),
    .B(_04213_),
    .CI(_04233_),
    .CO(_04234_),
    .S(_04235_));
 FA_X1 _09557_ (.A(_04236_),
    .B(\genblk1.gen_int_accumulation.int_adder.int_short_converted[10] ),
    .CI(\genblk1.gen_int_accumulation.int_adder.int_long_i[22] ),
    .CO(_04237_),
    .S(_04238_));
 FA_X1 _09558_ (.A(_04239_),
    .B(_04213_),
    .CI(_04240_),
    .CO(_04241_),
    .S(_04242_));
 FA_X1 _09559_ (.A(_04243_),
    .B(\genblk1.gen_int_accumulation.int_adder.int_short_converted[10] ),
    .CI(\genblk1.gen_int_accumulation.int_adder.int_long_i[26] ),
    .CO(_04244_),
    .S(_04245_));
 FA_X1 _09560_ (.A(_04246_),
    .B(\genblk1.gen_int_accumulation.int_adder.int_short_converted[10] ),
    .CI(\genblk1.gen_int_accumulation.int_adder.int_long_i[28] ),
    .CO(_04247_),
    .S(_04248_));
 FA_X1 _09561_ (.A(_04249_),
    .B(_04213_),
    .CI(_04250_),
    .CO(_04251_),
    .S(_04252_));
 HA_X1 _09562_ (.A(\genblk1.gen_int_accumulation.int_adder.int_short_converted[0] ),
    .B(\genblk1.gen_int_accumulation.int_adder.int_long_i[0] ),
    .CO(_04196_),
    .S(_04253_));
 HA_X1 _09563_ (.A(\genblk1.gen_int_accumulation.int_adder.int_short_converted[2] ),
    .B(\genblk1.gen_int_accumulation.int_adder.int_long_i[2] ),
    .CO(_04254_),
    .S(_04255_));
 HA_X1 _09564_ (.A(\genblk1.gen_int_accumulation.int_adder.int_short_converted[3] ),
    .B(\genblk1.gen_int_accumulation.int_adder.int_long_i[3] ),
    .CO(_04256_),
    .S(_04257_));
 HA_X1 _09565_ (.A(\genblk1.gen_int_accumulation.int_adder.int_short_converted[4] ),
    .B(\genblk1.gen_int_accumulation.int_adder.int_long_i[4] ),
    .CO(_04258_),
    .S(_04259_));
 HA_X1 _09566_ (.A(\genblk1.gen_int_accumulation.int_adder.int_short_converted[5] ),
    .B(\genblk1.gen_int_accumulation.int_adder.int_long_i[5] ),
    .CO(_04260_),
    .S(_04261_));
 HA_X1 _09567_ (.A(\genblk1.gen_int_accumulation.int_adder.int_short_converted[6] ),
    .B(\genblk1.gen_int_accumulation.int_adder.int_long_i[6] ),
    .CO(_04262_),
    .S(_04263_));
 HA_X1 _09568_ (.A(\genblk1.gen_int_accumulation.int_adder.int_short_converted[10] ),
    .B(\genblk1.gen_int_accumulation.int_adder.int_long_i[7] ),
    .CO(_04264_),
    .S(_04265_));
 HA_X1 _09569_ (.A(\genblk1.gen_int_accumulation.int_adder.int_short_converted[10] ),
    .B(\genblk1.gen_int_accumulation.int_adder.int_long_i[8] ),
    .CO(_04266_),
    .S(_04267_));
 HA_X1 _09570_ (.A(\genblk1.gen_int_accumulation.int_adder.int_short_converted[10] ),
    .B(\genblk1.gen_int_accumulation.int_adder.int_long_i[9] ),
    .CO(_04268_),
    .S(_04269_));
 HA_X1 _09571_ (.A(\genblk1.gen_int_accumulation.int_adder.int_short_converted[10] ),
    .B(\genblk1.gen_int_accumulation.int_adder.int_long_i[10] ),
    .CO(_04270_),
    .S(_04271_));
 HA_X1 _09572_ (.A(\genblk1.gen_int_accumulation.int_adder.int_short_converted[10] ),
    .B(\genblk1.gen_int_accumulation.int_adder.int_long_i[11] ),
    .CO(_04272_),
    .S(_04273_));
 HA_X1 _09573_ (.A(\genblk1.gen_int_accumulation.int_adder.int_short_converted[10] ),
    .B(\genblk1.gen_int_accumulation.int_adder.int_long_i[12] ),
    .CO(_04274_),
    .S(_04275_));
 HA_X1 _09574_ (.A(\genblk1.gen_int_accumulation.int_adder.int_short_converted[10] ),
    .B(\genblk1.gen_int_accumulation.int_adder.int_long_i[13] ),
    .CO(_04276_),
    .S(_04277_));
 HA_X1 _09575_ (.A(\genblk1.gen_int_accumulation.int_adder.int_short_converted[10] ),
    .B(\genblk1.gen_int_accumulation.int_adder.int_long_i[14] ),
    .CO(_04278_),
    .S(_04279_));
 HA_X1 _09576_ (.A(\genblk1.gen_int_accumulation.int_adder.int_short_converted[10] ),
    .B(\genblk1.gen_int_accumulation.int_adder.int_long_i[15] ),
    .CO(_04280_),
    .S(_04281_));
 HA_X1 _09577_ (.A(\genblk1.gen_int_accumulation.int_adder.int_short_converted[10] ),
    .B(\genblk1.gen_int_accumulation.int_adder.int_long_i[16] ),
    .CO(_04282_),
    .S(_04283_));
 HA_X1 _09578_ (.A(\genblk1.gen_int_accumulation.int_adder.int_short_converted[10] ),
    .B(\genblk1.gen_int_accumulation.int_adder.int_long_i[17] ),
    .CO(_04284_),
    .S(_04285_));
 HA_X1 _09579_ (.A(\genblk1.gen_int_accumulation.int_adder.int_short_converted[10] ),
    .B(\genblk1.gen_int_accumulation.int_adder.int_long_i[18] ),
    .CO(_04286_),
    .S(_04287_));
 HA_X1 _09580_ (.A(\genblk1.gen_int_accumulation.int_adder.int_short_converted[10] ),
    .B(\genblk1.gen_int_accumulation.int_adder.int_long_i[19] ),
    .CO(_04288_),
    .S(_04289_));
 HA_X1 _09581_ (.A(\genblk1.gen_int_accumulation.int_adder.int_short_converted[10] ),
    .B(\genblk1.gen_int_accumulation.int_adder.int_long_i[20] ),
    .CO(_04290_),
    .S(_04291_));
 HA_X1 _09582_ (.A(\genblk1.gen_int_accumulation.int_adder.int_short_converted[10] ),
    .B(\genblk1.gen_int_accumulation.int_adder.int_long_i[21] ),
    .CO(_04292_),
    .S(_04293_));
 HA_X1 _09583_ (.A(\genblk1.gen_int_accumulation.int_adder.int_short_converted[10] ),
    .B(\genblk1.gen_int_accumulation.int_adder.int_long_i[22] ),
    .CO(_04294_),
    .S(_04295_));
 HA_X1 _09584_ (.A(\genblk1.gen_int_accumulation.int_adder.int_short_converted[10] ),
    .B(\genblk1.gen_int_accumulation.int_adder.int_long_i[23] ),
    .CO(_04296_),
    .S(_04297_));
 HA_X1 _09585_ (.A(\genblk1.gen_int_accumulation.int_adder.int_short_converted[10] ),
    .B(\genblk1.gen_int_accumulation.int_adder.int_long_i[24] ),
    .CO(_04298_),
    .S(_04299_));
 HA_X1 _09586_ (.A(\genblk1.gen_int_accumulation.int_adder.int_short_converted[10] ),
    .B(\genblk1.gen_int_accumulation.int_adder.int_long_i[25] ),
    .CO(_04300_),
    .S(_04301_));
 HA_X1 _09587_ (.A(\genblk1.gen_int_accumulation.int_adder.int_short_converted[10] ),
    .B(\genblk1.gen_int_accumulation.int_adder.int_long_i[26] ),
    .CO(_04302_),
    .S(_04303_));
 HA_X1 _09588_ (.A(\genblk1.gen_int_accumulation.int_adder.int_short_converted[10] ),
    .B(\genblk1.gen_int_accumulation.int_adder.int_long_i[27] ),
    .CO(_04304_),
    .S(_04305_));
 HA_X1 _09589_ (.A(\genblk1.gen_int_accumulation.int_adder.int_short_converted[10] ),
    .B(\genblk1.gen_int_accumulation.int_adder.int_long_i[28] ),
    .CO(_04306_),
    .S(_04307_));
 HA_X1 _09590_ (.A(\genblk1.gen_int_accumulation.int_adder.int_short_converted[10] ),
    .B(\genblk1.gen_int_accumulation.int_adder.int_long_i[29] ),
    .CO(_04308_),
    .S(_04309_));
 DFFR_X1 _09591_ (.D(_00000_),
    .RN(net11),
    .CK(clknet_level_8_1_3434_clk_i),
    .Q(net30),
    .QN(_04160_));
 DFFR_X1 _09592_ (.D(_00001_),
    .RN(net11),
    .CK(clknet_level_8_1_3434_clk_i),
    .Q(net41),
    .QN(_04159_));
 DFFR_X1 _09593_ (.D(_00002_),
    .RN(net11),
    .CK(clknet_level_8_1_3434_clk_i),
    .Q(net52),
    .QN(_04158_));
 DFFR_X1 _09594_ (.D(_00003_),
    .RN(net11),
    .CK(clknet_level_8_1_3434_clk_i),
    .Q(net55),
    .QN(_04157_));
 DFFR_X1 _09595_ (.D(_00004_),
    .RN(net11),
    .CK(clknet_level_8_1_3434_clk_i),
    .Q(net56),
    .QN(_04156_));
 DFFR_X1 _09596_ (.D(_00005_),
    .RN(net11),
    .CK(clknet_level_8_1_4443_clk_i),
    .Q(net57),
    .QN(_04155_));
 DFFR_X1 _09597_ (.D(_00006_),
    .RN(net11),
    .CK(clknet_level_8_1_4443_clk_i),
    .Q(net58),
    .QN(_04154_));
 DFFR_X1 _09598_ (.D(_00007_),
    .RN(net11),
    .CK(clknet_level_8_1_4443_clk_i),
    .Q(net59),
    .QN(_04153_));
 DFFR_X1 _09599_ (.D(_00008_),
    .RN(net11),
    .CK(clknet_level_8_1_3434_clk_i),
    .Q(net60),
    .QN(_04152_));
 DFFR_X1 _09600_ (.D(_00009_),
    .RN(net11),
    .CK(clknet_level_8_1_4443_clk_i),
    .Q(net61),
    .QN(_04151_));
 DFFR_X1 _09601_ (.D(_00010_),
    .RN(net11),
    .CK(clknet_level_8_1_4443_clk_i),
    .Q(net31),
    .QN(_04150_));
 DFFR_X1 _09602_ (.D(_00011_),
    .RN(net11),
    .CK(clknet_level_8_1_4443_clk_i),
    .Q(net32),
    .QN(_04149_));
 DFFR_X1 _09603_ (.D(_00012_),
    .RN(net11),
    .CK(clknet_level_8_1_5452_clk_i),
    .Q(net33),
    .QN(_04148_));
 DFFR_X1 _09604_ (.D(_00013_),
    .RN(net11),
    .CK(clknet_level_8_1_6461_clk_i),
    .Q(net34),
    .QN(_04147_));
 DFFR_X1 _09605_ (.D(_00014_),
    .RN(net11),
    .CK(clknet_level_8_1_8479_clk_i),
    .Q(net35),
    .QN(_04146_));
 DFFR_X1 _09606_ (.D(_00015_),
    .RN(net11),
    .CK(clknet_level_8_1_8479_clk_i),
    .Q(net36),
    .QN(_04145_));
 DFFR_X1 _09607_ (.D(_00016_),
    .RN(net11),
    .CK(clknet_level_8_1_5452_clk_i),
    .Q(net37),
    .QN(_04144_));
 DFFR_X1 _09608_ (.D(_00017_),
    .RN(net11),
    .CK(clknet_level_8_1_5452_clk_i),
    .Q(net38),
    .QN(_04143_));
 DFFR_X1 _09609_ (.D(_00018_),
    .RN(net11),
    .CK(clknet_level_8_1_3434_clk_i),
    .Q(net39),
    .QN(_04142_));
 DFFR_X1 _09610_ (.D(_00019_),
    .RN(net11),
    .CK(clknet_level_8_1_3434_clk_i),
    .Q(net40),
    .QN(_04141_));
 DFFR_X1 _09611_ (.D(_00020_),
    .RN(net11),
    .CK(clknet_level_8_1_3434_clk_i),
    .Q(net42),
    .QN(_04140_));
 DFFR_X1 _09612_ (.D(_00021_),
    .RN(net11),
    .CK(clknet_level_8_1_3434_clk_i),
    .Q(net43),
    .QN(_04139_));
 DFFR_X1 _09613_ (.D(_00022_),
    .RN(net11),
    .CK(clknet_level_8_1_5452_clk_i),
    .Q(net44),
    .QN(_04138_));
 DFFR_X1 _09614_ (.D(_00023_),
    .RN(net11),
    .CK(clknet_level_8_1_5452_clk_i),
    .Q(net45),
    .QN(_04137_));
 DFFR_X1 _09615_ (.D(_00024_),
    .RN(net11),
    .CK(clknet_level_8_1_5452_clk_i),
    .Q(net46),
    .QN(_04136_));
 DFFR_X1 _09616_ (.D(_00025_),
    .RN(net11),
    .CK(clknet_level_8_1_7470_clk_i),
    .Q(net47),
    .QN(_04135_));
 DFFR_X1 _09617_ (.D(_00026_),
    .RN(net11),
    .CK(clknet_level_8_1_7470_clk_i),
    .Q(net48),
    .QN(_04134_));
 DFFR_X1 _09618_ (.D(_00027_),
    .RN(net11),
    .CK(clknet_level_8_1_7470_clk_i),
    .Q(net49),
    .QN(_04133_));
 DFFR_X1 _09619_ (.D(_00028_),
    .RN(net11),
    .CK(clknet_level_8_1_6461_clk_i),
    .Q(net50),
    .QN(_04132_));
 DFFR_X1 _09620_ (.D(_00029_),
    .RN(net11),
    .CK(clknet_level_8_1_8479_clk_i),
    .Q(net51),
    .QN(_04131_));
 DFFR_X1 _09621_ (.D(_00030_),
    .RN(net11),
    .CK(clknet_level_8_1_8479_clk_i),
    .Q(net53),
    .QN(_04130_));
 DFFR_X1 _09622_ (.D(_00031_),
    .RN(net11),
    .CK(clknet_level_8_1_8479_clk_i),
    .Q(net54),
    .QN(_04129_));
 DFFR_X2 _09623_ (.D(_00032_),
    .RN(net11),
    .CK(clknet_level_8_1_8479_clk_i),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[0] ),
    .QN(_04128_));
 DFFR_X2 _09624_ (.D(_00033_),
    .RN(net11),
    .CK(clknet_level_8_1_8479_clk_i),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[1] ),
    .QN(_04127_));
 DFFR_X2 _09625_ (.D(_00034_),
    .RN(net11),
    .CK(clknet_level_8_1_7470_clk_i),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[2] ),
    .QN(_04126_));
 DFFR_X2 _09626_ (.D(_00035_),
    .RN(net11),
    .CK(clknet_level_8_1_6461_clk_i),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[3] ),
    .QN(_04125_));
 DFFR_X2 _09627_ (.D(_00036_),
    .RN(net11),
    .CK(clknet_level_8_1_8479_clk_i),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[4] ),
    .QN(_04124_));
 DFFR_X2 _09628_ (.D(_00037_),
    .RN(net11),
    .CK(clknet_level_8_1_8479_clk_i),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[5] ),
    .QN(_04123_));
 DFFR_X2 _09629_ (.D(_00038_),
    .RN(net11),
    .CK(clknet_level_8_1_8479_clk_i),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[6] ),
    .QN(_04122_));
 DFFR_X2 _09630_ (.D(_00039_),
    .RN(net11),
    .CK(clknet_level_8_1_8479_clk_i),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[7] ),
    .QN(_04161_));
 DFFR_X1 _09631_ (.D(\rdata_o_n[0] ),
    .RN(net11),
    .CK(clknet_level_8_1_2425_clk_i),
    .Q(\genblk1.gen_int_accumulation.int_adder.int_short_converted[0] ),
    .QN(_04162_));
 DFFR_X1 _09632_ (.D(\rdata_o_n[1] ),
    .RN(net11),
    .CK(clknet_level_8_1_2425_clk_i),
    .Q(\genblk1.gen_int_accumulation.int_adder.int_short_converted[1] ),
    .QN(_04163_));
 DFFR_X1 _09633_ (.D(\rdata_o_n[2] ),
    .RN(net11),
    .CK(clknet_level_8_1_2425_clk_i),
    .Q(\genblk1.gen_int_accumulation.int_adder.int_short_converted[2] ),
    .QN(_04164_));
 DFFR_X1 _09634_ (.D(\rdata_o_n[3] ),
    .RN(net11),
    .CK(clknet_level_8_1_2425_clk_i),
    .Q(\genblk1.gen_int_accumulation.int_adder.int_short_converted[3] ),
    .QN(_04165_));
 DFFR_X1 _09635_ (.D(\rdata_o_n[4] ),
    .RN(net11),
    .CK(clknet_level_8_1_2425_clk_i),
    .Q(\genblk1.gen_int_accumulation.int_adder.int_short_converted[4] ),
    .QN(_04166_));
 DFFR_X1 _09636_ (.D(\rdata_o_n[5] ),
    .RN(net11),
    .CK(clknet_level_8_1_4443_clk_i),
    .Q(\genblk1.gen_int_accumulation.int_adder.int_short_converted[5] ),
    .QN(_04167_));
 DFFR_X1 _09637_ (.D(\rdata_o_n[6] ),
    .RN(net11),
    .CK(clknet_level_8_1_4443_clk_i),
    .Q(\genblk1.gen_int_accumulation.int_adder.int_short_converted[6] ),
    .QN(_04205_));
 DFFR_X2 _09638_ (.D(\rdata_o_n[7] ),
    .RN(net11),
    .CK(clknet_level_8_1_2425_clk_i),
    .Q(\genblk1.gen_int_accumulation.int_adder.int_short_converted[10] ),
    .QN(_04213_));
 DFFR_X1 _09639_ (.D(\result_int_n[0] ),
    .RN(net11),
    .CK(clknet_level_8_1_2425_clk_i),
    .Q(\genblk1.gen_int_accumulation.int_adder.int_long_i[0] ),
    .QN(_04168_));
 DFFR_X1 _09640_ (.D(\result_int_n[1] ),
    .RN(net11),
    .CK(clknet_level_8_1_4443_clk_i),
    .Q(\genblk1.gen_int_accumulation.int_adder.int_long_i[1] ),
    .QN(_04169_));
 DFFR_X1 _09641_ (.D(\result_int_n[2] ),
    .RN(net11),
    .CK(clknet_level_8_1_2425_clk_i),
    .Q(\genblk1.gen_int_accumulation.int_adder.int_long_i[2] ),
    .QN(_04170_));
 DFFR_X1 _09642_ (.D(\result_int_n[3] ),
    .RN(net11),
    .CK(clknet_level_8_1_2425_clk_i),
    .Q(\genblk1.gen_int_accumulation.int_adder.int_long_i[3] ),
    .QN(_04171_));
 DFFR_X1 _09643_ (.D(\result_int_n[4] ),
    .RN(net11),
    .CK(clknet_level_8_1_4443_clk_i),
    .Q(\genblk1.gen_int_accumulation.int_adder.int_long_i[4] ),
    .QN(_04172_));
 DFFR_X1 _09644_ (.D(\result_int_n[5] ),
    .RN(net11),
    .CK(clknet_level_8_1_2425_clk_i),
    .Q(\genblk1.gen_int_accumulation.int_adder.int_long_i[5] ),
    .QN(_04173_));
 DFFR_X1 _09645_ (.D(\result_int_n[6] ),
    .RN(net11),
    .CK(clknet_level_8_1_4443_clk_i),
    .Q(\genblk1.gen_int_accumulation.int_adder.int_long_i[6] ),
    .QN(_04206_));
 DFFR_X1 _09646_ (.D(\result_int_n[7] ),
    .RN(net11),
    .CK(clknet_level_8_1_4443_clk_i),
    .Q(\genblk1.gen_int_accumulation.int_adder.int_long_i[7] ),
    .QN(_04174_));
 DFFR_X1 _09647_ (.D(\result_int_n[8] ),
    .RN(net11),
    .CK(clknet_level_8_1_4443_clk_i),
    .Q(\genblk1.gen_int_accumulation.int_adder.int_long_i[8] ),
    .QN(_04175_));
 DFFR_X1 _09648_ (.D(\result_int_n[9] ),
    .RN(net11),
    .CK(clknet_level_8_1_4443_clk_i),
    .Q(\genblk1.gen_int_accumulation.int_adder.int_long_i[9] ),
    .QN(_04176_));
 DFFR_X1 _09649_ (.D(\result_int_n[10] ),
    .RN(net11),
    .CK(clknet_level_8_1_4443_clk_i),
    .Q(\genblk1.gen_int_accumulation.int_adder.int_long_i[10] ),
    .QN(_04214_));
 DFFR_X1 _09650_ (.D(\result_int_n[11] ),
    .RN(net11),
    .CK(clknet_level_8_1_4443_clk_i),
    .Q(\genblk1.gen_int_accumulation.int_adder.int_long_i[11] ),
    .QN(_04177_));
 DFFR_X1 _09651_ (.D(\result_int_n[12] ),
    .RN(net11),
    .CK(clknet_level_8_1_6461_clk_i),
    .Q(\genblk1.gen_int_accumulation.int_adder.int_long_i[12] ),
    .QN(_04218_));
 DFFR_X1 _09652_ (.D(\result_int_n[13] ),
    .RN(net11),
    .CK(clknet_level_8_1_7470_clk_i),
    .Q(\genblk1.gen_int_accumulation.int_adder.int_long_i[13] ),
    .QN(_04178_));
 DFFR_X1 _09653_ (.D(\result_int_n[14] ),
    .RN(net11),
    .CK(clknet_level_8_1_7470_clk_i),
    .Q(\genblk1.gen_int_accumulation.int_adder.int_long_i[14] ),
    .QN(_04222_));
 DFFR_X1 _09654_ (.D(\result_int_n[15] ),
    .RN(net11),
    .CK(clknet_level_8_1_7470_clk_i),
    .Q(\genblk1.gen_int_accumulation.int_adder.int_long_i[15] ),
    .QN(_04179_));
 DFFR_X1 _09655_ (.D(\result_int_n[16] ),
    .RN(net11),
    .CK(clknet_level_8_1_5452_clk_i),
    .Q(\genblk1.gen_int_accumulation.int_adder.int_long_i[16] ),
    .QN(_04180_));
 DFFR_X1 _09656_ (.D(\result_int_n[17] ),
    .RN(net11),
    .CK(clknet_level_8_1_5452_clk_i),
    .Q(\genblk1.gen_int_accumulation.int_adder.int_long_i[17] ),
    .QN(_04181_));
 DFFR_X1 _09657_ (.D(\result_int_n[18] ),
    .RN(net11),
    .CK(clknet_level_8_1_3434_clk_i),
    .Q(\genblk1.gen_int_accumulation.int_adder.int_long_i[18] ),
    .QN(_04229_));
 DFFR_X1 _09658_ (.D(\result_int_n[19] ),
    .RN(net11),
    .CK(clknet_level_8_1_3434_clk_i),
    .Q(\genblk1.gen_int_accumulation.int_adder.int_long_i[19] ),
    .QN(_04182_));
 DFFR_X1 _09659_ (.D(\result_int_n[20] ),
    .RN(net11),
    .CK(clknet_level_8_1_2425_clk_i),
    .Q(\genblk1.gen_int_accumulation.int_adder.int_long_i[20] ),
    .QN(_04233_));
 DFFR_X1 _09660_ (.D(\result_int_n[21] ),
    .RN(net11),
    .CK(clknet_level_8_1_2425_clk_i),
    .Q(\genblk1.gen_int_accumulation.int_adder.int_long_i[21] ),
    .QN(_04183_));
 DFFR_X1 _09661_ (.D(\result_int_n[22] ),
    .RN(net11),
    .CK(clknet_level_8_1_7470_clk_i),
    .Q(\genblk1.gen_int_accumulation.int_adder.int_long_i[22] ),
    .QN(_04184_));
 DFFR_X1 _09662_ (.D(\result_int_n[23] ),
    .RN(net11),
    .CK(clknet_level_8_1_7470_clk_i),
    .Q(\genblk1.gen_int_accumulation.int_adder.int_long_i[23] ),
    .QN(_04185_));
 DFFR_X1 _09663_ (.D(\result_int_n[24] ),
    .RN(net11),
    .CK(clknet_level_8_1_5452_clk_i),
    .Q(\genblk1.gen_int_accumulation.int_adder.int_long_i[24] ),
    .QN(_04240_));
 DFFR_X1 _09664_ (.D(\result_int_n[25] ),
    .RN(net11),
    .CK(clknet_level_8_1_7470_clk_i),
    .Q(\genblk1.gen_int_accumulation.int_adder.int_long_i[25] ),
    .QN(_04186_));
 DFFR_X1 _09665_ (.D(\result_int_n[26] ),
    .RN(net11),
    .CK(clknet_level_8_1_8479_clk_i),
    .Q(\genblk1.gen_int_accumulation.int_adder.int_long_i[26] ),
    .QN(_04187_));
 DFFR_X1 _09666_ (.D(\result_int_n[27] ),
    .RN(net11),
    .CK(clknet_level_8_1_8479_clk_i),
    .Q(\genblk1.gen_int_accumulation.int_adder.int_long_i[27] ),
    .QN(_04188_));
 DFFR_X1 _09667_ (.D(\result_int_n[28] ),
    .RN(net11),
    .CK(clknet_level_8_1_6461_clk_i),
    .Q(\genblk1.gen_int_accumulation.int_adder.int_long_i[28] ),
    .QN(_04189_));
 DFFR_X1 _09668_ (.D(\result_int_n[29] ),
    .RN(net11),
    .CK(clknet_level_8_1_6461_clk_i),
    .Q(\genblk1.gen_int_accumulation.int_adder.int_long_i[29] ),
    .QN(_04190_));
 DFFR_X1 _09669_ (.D(\result_int_n[30] ),
    .RN(net11),
    .CK(clknet_level_8_1_6461_clk_i),
    .Q(\genblk1.gen_int_accumulation.int_adder.int_long_i[30] ),
    .QN(_04250_));
 DFFR_X1 _09670_ (.D(\result_int_n[31] ),
    .RN(net11),
    .CK(clknet_level_8_1_8479_clk_i),
    .Q(\genblk1.gen_int_accumulation.int_adder.int_long_i[31] ),
    .QN(_04121_));
 DFFR_X2 _09671_ (.D(_00040_),
    .RN(net11),
    .CK(clknet_level_8_1_18_clk_i),
    .Q(net62),
    .QN(_04191_));
 DFFR_X1 _09672_ (.D(\caddr_n[0] ),
    .RN(net11),
    .CK(clknet_level_8_1_18_clk_i),
    .Q(\caddr_q[0] ),
    .QN(_04192_));
 DFFR_X1 _09673_ (.D(\caddr_n[1] ),
    .RN(net11),
    .CK(clknet_level_8_1_18_clk_i),
    .Q(\caddr_q[1] ),
    .QN(_04193_));
 DFFR_X1 _09674_ (.D(\caddr_n[2] ),
    .RN(net11),
    .CK(clknet_level_8_1_18_clk_i),
    .Q(\caddr_q[2] ),
    .QN(_04194_));
 DFFR_X1 _09675_ (.D(\caddr_n[3] ),
    .RN(net11),
    .CK(clknet_level_8_1_18_clk_i),
    .Q(\caddr_q[3] ),
    .QN(_04195_));
 DFFR_X1 _09676_ (.D(\caddr_n[4] ),
    .RN(net11),
    .CK(clknet_level_8_1_18_clk_i),
    .Q(\caddr_q[4] ),
    .QN(_04120_));
 DLH_X1 _09677_ (.D(net321),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[13][0] ));
 DLH_X1 _09678_ (.D(net310),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[13][1] ));
 DLH_X1 _09679_ (.D(net308),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[13][2] ));
 DLH_X1 _09680_ (.D(net302),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[13][3] ));
 DLH_X1 _09681_ (.D(net293),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[13][4] ));
 DLH_X1 _09682_ (.D(net291),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[13][5] ));
 DLH_X1 _09683_ (.D(net283),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[13][6] ));
 DLH_X1 _09684_ (.D(net275),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[13][7] ));
 DLH_X1 _09685_ (.D(net321),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[1][0] ));
 DLH_X1 _09686_ (.D(net310),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[1][1] ));
 DLH_X1 _09687_ (.D(net308),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[1][2] ));
 DLH_X1 _09688_ (.D(net302),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[1][3] ));
 DLH_X1 _09689_ (.D(net293),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[1][4] ));
 DLH_X1 _09690_ (.D(net291),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[1][5] ));
 DLH_X1 _09691_ (.D(net283),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[1][6] ));
 DLH_X1 _09692_ (.D(net275),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[1][7] ));
 DLH_X1 _09693_ (.D(net321),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[26][0] ));
 DLH_X1 _09694_ (.D(net310),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[26][1] ));
 DLH_X1 _09695_ (.D(net308),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[26][2] ));
 DLH_X1 _09696_ (.D(net302),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[26][3] ));
 DLH_X1 _09697_ (.D(net293),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[26][4] ));
 DLH_X1 _09698_ (.D(net291),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[26][5] ));
 DLH_X1 _09699_ (.D(net283),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[26][6] ));
 DLH_X1 _09700_ (.D(net275),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[26][7] ));
 DLH_X1 _09701_ (.D(net321),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[9][0] ));
 DLH_X1 _09702_ (.D(net310),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[9][1] ));
 DLH_X1 _09703_ (.D(net308),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[9][2] ));
 DLH_X1 _09704_ (.D(net302),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[9][3] ));
 DLH_X1 _09705_ (.D(net293),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[9][4] ));
 DLH_X1 _09706_ (.D(net291),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[9][5] ));
 DLH_X1 _09707_ (.D(net283),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[9][6] ));
 DLH_X1 _09708_ (.D(net275),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[9][7] ));
 DLH_X1 _09709_ (.D(net320),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[0][0] ));
 DLH_X1 _09710_ (.D(net311),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[0][1] ));
 DLH_X1 _09711_ (.D(net305),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[0][2] ));
 DLH_X1 _09712_ (.D(net300),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[0][3] ));
 DLH_X1 _09713_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[4] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[0][4] ));
 DLH_X1 _09714_ (.D(net292),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[0][5] ));
 DLH_X1 _09715_ (.D(net285),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[0][6] ));
 DLH_X1 _09716_ (.D(net275),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[0][7] ));
 DLH_X1 _09717_ (.D(net321),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[20][0] ));
 DLH_X1 _09718_ (.D(net310),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[20][1] ));
 DLH_X1 _09719_ (.D(net308),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[20][2] ));
 DLH_X1 _09720_ (.D(net302),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[20][3] ));
 DLH_X1 _09721_ (.D(net293),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[20][4] ));
 DLH_X1 _09722_ (.D(net291),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[20][5] ));
 DLH_X1 _09723_ (.D(net283),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[20][6] ));
 DLH_X1 _09724_ (.D(net275),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[20][7] ));
 DLH_X1 _09725_ (.D(net321),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[2][0] ));
 DLH_X1 _09726_ (.D(net310),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[2][1] ));
 DLH_X1 _09727_ (.D(net308),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[2][2] ));
 DLH_X1 _09728_ (.D(net302),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[2][3] ));
 DLH_X1 _09729_ (.D(net293),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[2][4] ));
 DLH_X1 _09730_ (.D(net291),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[2][5] ));
 DLH_X1 _09731_ (.D(net283),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[2][6] ));
 DLH_X1 _09732_ (.D(net275),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[2][7] ));
 DLH_X1 _09733_ (.D(net321),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[25][0] ));
 DLH_X1 _09734_ (.D(net310),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[25][1] ));
 DLH_X1 _09735_ (.D(net308),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[25][2] ));
 DLH_X1 _09736_ (.D(net302),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[25][3] ));
 DLH_X1 _09737_ (.D(net293),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[25][4] ));
 DLH_X1 _09738_ (.D(net291),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[25][5] ));
 DLH_X1 _09739_ (.D(net283),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[25][6] ));
 DLH_X1 _09740_ (.D(net275),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[25][7] ));
 DLH_X1 _09741_ (.D(net321),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[10][0] ));
 DLH_X1 _09742_ (.D(net310),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[10][1] ));
 DLH_X1 _09743_ (.D(net308),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[10][2] ));
 DLH_X1 _09744_ (.D(net302),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[10][3] ));
 DLH_X1 _09745_ (.D(net293),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[10][4] ));
 DLH_X1 _09746_ (.D(net291),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[10][5] ));
 DLH_X1 _09747_ (.D(net283),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[10][6] ));
 DLH_X1 _09748_ (.D(net275),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[10][7] ));
 DLH_X1 _09749_ (.D(net321),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[3][0] ));
 DLH_X1 _09750_ (.D(net310),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[3][1] ));
 DLH_X1 _09751_ (.D(net308),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[3][2] ));
 DLH_X1 _09752_ (.D(net302),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[3][3] ));
 DLH_X1 _09753_ (.D(net293),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[3][4] ));
 DLH_X1 _09754_ (.D(net291),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[3][5] ));
 DLH_X1 _09755_ (.D(net283),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[3][6] ));
 DLH_X1 _09756_ (.D(net275),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[3][7] ));
 DLH_X1 _09757_ (.D(net321),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[16][0] ));
 DLH_X1 _09758_ (.D(net310),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[16][1] ));
 DLH_X1 _09759_ (.D(net308),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[16][2] ));
 DLH_X1 _09760_ (.D(net302),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[16][3] ));
 DLH_X1 _09761_ (.D(net293),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[16][4] ));
 DLH_X1 _09762_ (.D(net291),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[16][5] ));
 DLH_X1 _09763_ (.D(net283),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[16][6] ));
 DLH_X1 _09764_ (.D(net275),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[16][7] ));
 DLH_X1 _09765_ (.D(net321),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[24][0] ));
 DLH_X1 _09766_ (.D(net310),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[24][1] ));
 DLH_X1 _09767_ (.D(net308),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[24][2] ));
 DLH_X1 _09768_ (.D(net302),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[24][3] ));
 DLH_X1 _09769_ (.D(net293),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[24][4] ));
 DLH_X1 _09770_ (.D(net291),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[24][5] ));
 DLH_X1 _09771_ (.D(net283),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[24][6] ));
 DLH_X1 _09772_ (.D(net275),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[24][7] ));
 DLH_X1 _09773_ (.D(net321),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[4][0] ));
 DLH_X1 _09774_ (.D(net310),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[4][1] ));
 DLH_X1 _09775_ (.D(net308),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[4][2] ));
 DLH_X1 _09776_ (.D(net302),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[4][3] ));
 DLH_X1 _09777_ (.D(net293),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[4][4] ));
 DLH_X1 _09778_ (.D(net291),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[4][5] ));
 DLH_X1 _09779_ (.D(net283),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[4][6] ));
 DLH_X1 _09780_ (.D(net275),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[4][7] ));
 DLH_X1 _09781_ (.D(net321),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[15][0] ));
 DLH_X1 _09782_ (.D(net310),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[15][1] ));
 DLH_X1 _09783_ (.D(net308),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[15][2] ));
 DLH_X1 _09784_ (.D(net302),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[15][3] ));
 DLH_X1 _09785_ (.D(net293),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[15][4] ));
 DLH_X1 _09786_ (.D(net291),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[15][5] ));
 DLH_X1 _09787_ (.D(net283),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[15][6] ));
 DLH_X1 _09788_ (.D(net275),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[15][7] ));
 DLH_X1 _09789_ (.D(net321),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[11][0] ));
 DLH_X1 _09790_ (.D(net310),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[11][1] ));
 DLH_X1 _09791_ (.D(net308),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[11][2] ));
 DLH_X1 _09792_ (.D(net302),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[11][3] ));
 DLH_X1 _09793_ (.D(net293),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[11][4] ));
 DLH_X1 _09794_ (.D(net291),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[11][5] ));
 DLH_X1 _09795_ (.D(net283),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[11][6] ));
 DLH_X1 _09796_ (.D(net275),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[11][7] ));
 DLH_X1 _09797_ (.D(net321),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[5][0] ));
 DLH_X1 _09798_ (.D(net310),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[5][1] ));
 DLH_X1 _09799_ (.D(net308),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[5][2] ));
 DLH_X1 _09800_ (.D(net302),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[5][3] ));
 DLH_X1 _09801_ (.D(net293),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[5][4] ));
 DLH_X1 _09802_ (.D(net291),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[5][5] ));
 DLH_X1 _09803_ (.D(net283),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[5][6] ));
 DLH_X1 _09804_ (.D(net275),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[5][7] ));
 DLH_X1 _09805_ (.D(net321),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[23][0] ));
 DLH_X1 _09806_ (.D(net310),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[23][1] ));
 DLH_X1 _09807_ (.D(net308),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[23][2] ));
 DLH_X1 _09808_ (.D(net302),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[23][3] ));
 DLH_X1 _09809_ (.D(net293),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[23][4] ));
 DLH_X1 _09810_ (.D(net291),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[23][5] ));
 DLH_X1 _09811_ (.D(net283),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[23][6] ));
 DLH_X1 _09812_ (.D(net275),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[23][7] ));
 DLH_X1 _09813_ (.D(net321),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[19][0] ));
 DLH_X1 _09814_ (.D(net310),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[19][1] ));
 DLH_X1 _09815_ (.D(net308),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[19][2] ));
 DLH_X1 _09816_ (.D(net302),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[19][3] ));
 DLH_X1 _09817_ (.D(net293),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[19][4] ));
 DLH_X1 _09818_ (.D(net291),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[19][5] ));
 DLH_X1 _09819_ (.D(net283),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[19][6] ));
 DLH_X1 _09820_ (.D(net275),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[19][7] ));
 DLH_X1 _09821_ (.D(net321),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[31][0] ));
 DLH_X1 _09822_ (.D(net310),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[31][1] ));
 DLH_X1 _09823_ (.D(net308),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[31][2] ));
 DLH_X1 _09824_ (.D(net302),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[31][3] ));
 DLH_X1 _09825_ (.D(net293),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[31][4] ));
 DLH_X1 _09826_ (.D(net291),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[31][5] ));
 DLH_X1 _09827_ (.D(net283),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[31][6] ));
 DLH_X1 _09828_ (.D(net275),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[31][7] ));
 DLH_X1 _09829_ (.D(net321),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[6][0] ));
 DLH_X1 _09830_ (.D(net310),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[6][1] ));
 DLH_X1 _09831_ (.D(net308),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[6][2] ));
 DLH_X1 _09832_ (.D(net302),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[6][3] ));
 DLH_X1 _09833_ (.D(net293),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[6][4] ));
 DLH_X1 _09834_ (.D(net291),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[6][5] ));
 DLH_X1 _09835_ (.D(net283),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[6][6] ));
 DLH_X1 _09836_ (.D(net275),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[6][7] ));
 DLH_X1 _09837_ (.D(net321),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[14][0] ));
 DLH_X1 _09838_ (.D(net310),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[14][1] ));
 DLH_X1 _09839_ (.D(net308),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[14][2] ));
 DLH_X1 _09840_ (.D(net302),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[14][3] ));
 DLH_X1 _09841_ (.D(net293),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[14][4] ));
 DLH_X1 _09842_ (.D(net291),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[14][5] ));
 DLH_X1 _09843_ (.D(net283),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[14][6] ));
 DLH_X1 _09844_ (.D(net275),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[14][7] ));
 DLH_X1 _09845_ (.D(net321),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[30][0] ));
 DLH_X1 _09846_ (.D(net310),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[30][1] ));
 DLH_X1 _09847_ (.D(net308),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[30][2] ));
 DLH_X1 _09848_ (.D(net302),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[30][3] ));
 DLH_X1 _09849_ (.D(net293),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[30][4] ));
 DLH_X1 _09850_ (.D(net291),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[30][5] ));
 DLH_X1 _09851_ (.D(net283),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[30][6] ));
 DLH_X1 _09852_ (.D(net275),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[30][7] ));
 DLH_X1 _09853_ (.D(net321),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[22][0] ));
 DLH_X1 _09854_ (.D(net310),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[22][1] ));
 DLH_X1 _09855_ (.D(net308),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[22][2] ));
 DLH_X1 _09856_ (.D(net302),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[22][3] ));
 DLH_X1 _09857_ (.D(net293),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[22][4] ));
 DLH_X1 _09858_ (.D(net291),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[22][5] ));
 DLH_X1 _09859_ (.D(net283),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[22][6] ));
 DLH_X1 _09860_ (.D(net275),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[22][7] ));
 DLH_X1 _09861_ (.D(net321),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[7][0] ));
 DLH_X1 _09862_ (.D(net310),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[7][1] ));
 DLH_X1 _09863_ (.D(net308),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[7][2] ));
 DLH_X1 _09864_ (.D(net302),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[7][3] ));
 DLH_X1 _09865_ (.D(net293),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[7][4] ));
 DLH_X1 _09866_ (.D(net291),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[7][5] ));
 DLH_X1 _09867_ (.D(net283),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[7][6] ));
 DLH_X1 _09868_ (.D(net275),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[7][7] ));
 DLH_X1 _09869_ (.D(net321),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[29][0] ));
 DLH_X1 _09870_ (.D(net310),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[29][1] ));
 DLH_X1 _09871_ (.D(net308),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[29][2] ));
 DLH_X1 _09872_ (.D(net302),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[29][3] ));
 DLH_X1 _09873_ (.D(net293),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[29][4] ));
 DLH_X1 _09874_ (.D(net291),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[29][5] ));
 DLH_X1 _09875_ (.D(net283),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[29][6] ));
 DLH_X1 _09876_ (.D(net275),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[29][7] ));
 DLH_X1 _09877_ (.D(net321),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[12][0] ));
 DLH_X1 _09878_ (.D(net310),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[12][1] ));
 DLH_X1 _09879_ (.D(net308),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[12][2] ));
 DLH_X1 _09880_ (.D(net302),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[12][3] ));
 DLH_X1 _09881_ (.D(net293),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[12][4] ));
 DLH_X1 _09882_ (.D(net291),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[12][5] ));
 DLH_X1 _09883_ (.D(net283),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[12][6] ));
 DLH_X1 _09884_ (.D(net275),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[12][7] ));
 DLH_X1 _09885_ (.D(net321),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[17][0] ));
 DLH_X1 _09886_ (.D(net310),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[17][1] ));
 DLH_X1 _09887_ (.D(net308),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[17][2] ));
 DLH_X1 _09888_ (.D(net302),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[17][3] ));
 DLH_X1 _09889_ (.D(net293),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[17][4] ));
 DLH_X1 _09890_ (.D(net291),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[17][5] ));
 DLH_X1 _09891_ (.D(net283),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[17][6] ));
 DLH_X1 _09892_ (.D(net275),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[17][7] ));
 DLH_X1 _09893_ (.D(net321),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[28][0] ));
 DLH_X1 _09894_ (.D(net310),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[28][1] ));
 DLH_X1 _09895_ (.D(net308),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[28][2] ));
 DLH_X1 _09896_ (.D(net302),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[28][3] ));
 DLH_X1 _09897_ (.D(net293),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[28][4] ));
 DLH_X1 _09898_ (.D(net291),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[28][5] ));
 DLH_X1 _09899_ (.D(net283),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[28][6] ));
 DLH_X1 _09900_ (.D(net275),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[28][7] ));
 DLH_X1 _09901_ (.D(net321),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[8][0] ));
 DLH_X1 _09902_ (.D(net310),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[8][1] ));
 DLH_X1 _09903_ (.D(net308),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[8][2] ));
 DLH_X1 _09904_ (.D(net302),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[8][3] ));
 DLH_X1 _09905_ (.D(net293),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[8][4] ));
 DLH_X1 _09906_ (.D(net291),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[8][5] ));
 DLH_X1 _09907_ (.D(net283),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[8][6] ));
 DLH_X1 _09908_ (.D(net275),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[8][7] ));
 DLH_X1 _09909_ (.D(net321),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[21][0] ));
 DLH_X1 _09910_ (.D(net310),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[21][1] ));
 DLH_X1 _09911_ (.D(net308),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[21][2] ));
 DLH_X1 _09912_ (.D(net302),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[21][3] ));
 DLH_X1 _09913_ (.D(net293),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[21][4] ));
 DLH_X1 _09914_ (.D(net291),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[21][5] ));
 DLH_X1 _09915_ (.D(net283),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[21][6] ));
 DLH_X1 _09916_ (.D(net275),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[21][7] ));
 DLH_X1 _09917_ (.D(net321),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[27][0] ));
 DLH_X1 _09918_ (.D(net310),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[27][1] ));
 DLH_X1 _09919_ (.D(net308),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[27][2] ));
 DLH_X1 _09920_ (.D(net302),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[27][3] ));
 DLH_X1 _09921_ (.D(net293),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[27][4] ));
 DLH_X1 _09922_ (.D(net291),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[27][5] ));
 DLH_X1 _09923_ (.D(net283),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[27][6] ));
 DLH_X1 _09924_ (.D(net275),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[27][7] ));
 DLH_X1 _09925_ (.D(net321),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[18][0] ));
 DLH_X1 _09926_ (.D(net310),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[18][1] ));
 DLH_X1 _09927_ (.D(net308),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[18][2] ));
 DLH_X1 _09928_ (.D(net302),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[18][3] ));
 DLH_X1 _09929_ (.D(net293),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[18][4] ));
 DLH_X1 _09930_ (.D(net291),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[18][5] ));
 DLH_X1 _09931_ (.D(net283),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[18][6] ));
 DLH_X1 _09932_ (.D(net275),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.mem[18][7] ));
 DLL_X1 _09933_ (.D(\lut.gen_sub_units_scm.__15.sub_unit_i.cg_we_global.en_i ),
    .GN(clknet_level_5_1_3218__00532_),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.cg_we_global.clk_en ));
 DLL_X1 _09934_ (.D(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__0.cg_i.en_i ),
    .GN(clknet_level_2_1_6236__00534_),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_en ));
 DLL_X1 _09935_ (.D(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__1.cg_i.en_i ),
    .GN(clknet_level_2_1_1221__00534_),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_en ));
 DLL_X1 _09936_ (.D(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__2.cg_i.en_i ),
    .GN(clknet_level_2_1_4230__00534_),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_en ));
 DLL_X1 _09937_ (.D(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__3.cg_i.en_i ),
    .GN(clknet_level_2_1_2224__00534_),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_en ));
 DLL_X1 _09938_ (.D(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__4.cg_i.en_i ),
    .GN(clknet_level_2_1_2224__00534_),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_en ));
 DLL_X1 _09939_ (.D(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__5.cg_i.en_i ),
    .GN(clknet_level_2_1_4230__00534_),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_en ));
 DLL_X1 _09940_ (.D(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__6.cg_i.en_i ),
    .GN(clknet_level_2_1_6236__00534_),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_en ));
 DLL_X1 _09941_ (.D(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__7.cg_i.en_i ),
    .GN(clknet_level_2_1_4230__00534_),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_en ));
 DLL_X1 _09942_ (.D(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__8.cg_i.en_i ),
    .GN(clknet_level_2_1_2224__00534_),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_en ));
 DLL_X1 _09943_ (.D(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__9.cg_i.en_i ),
    .GN(clknet_level_2_1_7239__00534_),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_en ));
 DLL_X1 _09944_ (.D(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__10.cg_i.en_i ),
    .GN(clknet_level_2_1_5233__00534_),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_en ));
 DLL_X1 _09945_ (.D(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__11.cg_i.en_i ),
    .GN(clknet_level_2_1_8242__00534_),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_en ));
 DLL_X1 _09946_ (.D(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__12.cg_i.en_i ),
    .GN(clknet_level_2_1_3227__00534_),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_en ));
 DLL_X1 _09947_ (.D(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__13.cg_i.en_i ),
    .GN(clknet_level_2_1_1221__00534_),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_en ));
 DLL_X1 _09948_ (.D(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__14.cg_i.en_i ),
    .GN(clknet_level_2_1_3227__00534_),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_en ));
 DLL_X1 _09949_ (.D(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__15.cg_i.en_i ),
    .GN(clknet_level_2_1_3227__00534_),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_en ));
 DLL_X1 _09950_ (.D(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__16.cg_i.en_i ),
    .GN(clknet_level_2_1_1221__00534_),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_en ));
 DLL_X1 _09951_ (.D(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__17.cg_i.en_i ),
    .GN(clknet_level_2_1_7239__00534_),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_en ));
 DLL_X1 _09952_ (.D(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__18.cg_i.en_i ),
    .GN(clknet_level_2_1_1221__00534_),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_en ));
 DLL_X1 _09953_ (.D(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__19.cg_i.en_i ),
    .GN(clknet_level_2_1_3227__00534_),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_en ));
 DLL_X1 _09954_ (.D(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__20.cg_i.en_i ),
    .GN(clknet_level_2_1_4230__00534_),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_en ));
 DLL_X1 _09955_ (.D(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__21.cg_i.en_i ),
    .GN(clknet_level_2_1_8242__00534_),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_en ));
 DLL_X1 _09956_ (.D(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__22.cg_i.en_i ),
    .GN(clknet_level_2_1_3227__00534_),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_en ));
 DLL_X1 _09957_ (.D(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__23.cg_i.en_i ),
    .GN(clknet_level_2_1_5233__00534_),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_en ));
 DLL_X1 _09958_ (.D(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__24.cg_i.en_i ),
    .GN(clknet_level_2_1_2224__00534_),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_en ));
 DLL_X1 _09959_ (.D(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__25.cg_i.en_i ),
    .GN(clknet_level_2_1_6236__00534_),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_en ));
 DLL_X1 _09960_ (.D(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__26.cg_i.en_i ),
    .GN(clknet_level_2_1_2224__00534_),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_en ));
 DLL_X1 _09961_ (.D(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__27.cg_i.en_i ),
    .GN(clknet_level_2_1_6236__00534_),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_en ));
 DLL_X1 _09962_ (.D(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__28.cg_i.en_i ),
    .GN(clknet_level_2_1_8242__00534_),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_en ));
 DLL_X1 _09963_ (.D(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__29.cg_i.en_i ),
    .GN(clknet_level_2_1_8242__00534_),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_en ));
 DLL_X1 _09964_ (.D(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__30.cg_i.en_i ),
    .GN(clknet_level_2_1_4230__00534_),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_en ));
 DLL_X1 _09965_ (.D(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__31.cg_i.en_i ),
    .GN(clknet_level_2_1_5233__00534_),
    .Q(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_en ));
 DLH_X1 _09966_ (.D(net316),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[13][0] ));
 DLH_X1 _09967_ (.D(net313),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[13][1] ));
 DLH_X1 _09968_ (.D(net306),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[13][2] ));
 DLH_X1 _09969_ (.D(net298),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[13][3] ));
 DLH_X1 _09970_ (.D(net295),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[13][4] ));
 DLH_X1 _09971_ (.D(net288),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[13][5] ));
 DLH_X1 _09972_ (.D(net282),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[13][6] ));
 DLH_X1 _09973_ (.D(net276),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[13][7] ));
 DLH_X1 _09974_ (.D(net316),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[1][0] ));
 DLH_X1 _09975_ (.D(net313),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[1][1] ));
 DLH_X1 _09976_ (.D(net304),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[1][2] ));
 DLH_X1 _09977_ (.D(net303),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[1][3] ));
 DLH_X1 _09978_ (.D(net295),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[1][4] ));
 DLH_X1 _09979_ (.D(net288),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[1][5] ));
 DLH_X1 _09980_ (.D(net284),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[1][6] ));
 DLH_X1 _09981_ (.D(net277),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[1][7] ));
 DLH_X1 _09982_ (.D(net319),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[26][0] ));
 DLH_X1 _09983_ (.D(net313),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[26][1] ));
 DLH_X1 _09984_ (.D(net304),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[26][2] ));
 DLH_X1 _09985_ (.D(net298),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[26][3] ));
 DLH_X1 _09986_ (.D(net295),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[26][4] ));
 DLH_X1 _09987_ (.D(net292),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[26][5] ));
 DLH_X1 _09988_ (.D(net284),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[26][6] ));
 DLH_X1 _09989_ (.D(net276),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[26][7] ));
 DLH_X1 _09990_ (.D(net316),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[9][0] ));
 DLH_X1 _09991_ (.D(net313),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[9][1] ));
 DLH_X1 _09992_ (.D(net304),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[9][2] ));
 DLH_X1 _09993_ (.D(net298),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[9][3] ));
 DLH_X1 _09994_ (.D(net295),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[9][4] ));
 DLH_X1 _09995_ (.D(net288),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[9][5] ));
 DLH_X1 _09996_ (.D(net282),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[9][6] ));
 DLH_X1 _09997_ (.D(net279),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[9][7] ));
 DLH_X1 _09998_ (.D(net316),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[0][0] ));
 DLH_X1 _09999_ (.D(net311),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[0][1] ));
 DLH_X1 _10000_ (.D(net306),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[0][2] ));
 DLH_X1 _10001_ (.D(net303),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[0][3] ));
 DLH_X1 _10002_ (.D(net295),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[0][4] ));
 DLH_X1 _10003_ (.D(net288),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[0][5] ));
 DLH_X1 _10004_ (.D(net284),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[0][6] ));
 DLH_X1 _10005_ (.D(net277),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[0][7] ));
 DLH_X1 _10006_ (.D(net319),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[20][0] ));
 DLH_X1 _10007_ (.D(net313),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[20][1] ));
 DLH_X1 _10008_ (.D(net306),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[20][2] ));
 DLH_X1 _10009_ (.D(net298),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[20][3] ));
 DLH_X1 _10010_ (.D(net295),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[20][4] ));
 DLH_X1 _10011_ (.D(net288),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[20][5] ));
 DLH_X1 _10012_ (.D(net284),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[20][6] ));
 DLH_X1 _10013_ (.D(net277),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[20][7] ));
 DLH_X1 _10014_ (.D(net316),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[2][0] ));
 DLH_X1 _10015_ (.D(net313),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[2][1] ));
 DLH_X1 _10016_ (.D(net306),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[2][2] ));
 DLH_X1 _10017_ (.D(net298),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[2][3] ));
 DLH_X1 _10018_ (.D(net295),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[2][4] ));
 DLH_X1 _10019_ (.D(net288),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[2][5] ));
 DLH_X1 _10020_ (.D(net284),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[2][6] ));
 DLH_X1 _10021_ (.D(net276),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[2][7] ));
 DLH_X1 _10022_ (.D(net319),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[25][0] ));
 DLH_X1 _10023_ (.D(net313),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[25][1] ));
 DLH_X1 _10024_ (.D(net306),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[25][2] ));
 DLH_X1 _10025_ (.D(net298),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[25][3] ));
 DLH_X1 _10026_ (.D(net295),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[25][4] ));
 DLH_X1 _10027_ (.D(net288),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[25][5] ));
 DLH_X1 _10028_ (.D(net284),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[25][6] ));
 DLH_X1 _10029_ (.D(net276),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[25][7] ));
 DLH_X1 _10030_ (.D(net319),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[10][0] ));
 DLH_X1 _10031_ (.D(net313),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[10][1] ));
 DLH_X1 _10032_ (.D(net304),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[10][2] ));
 DLH_X1 _10033_ (.D(net298),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[10][3] ));
 DLH_X1 _10034_ (.D(net295),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[10][4] ));
 DLH_X1 _10035_ (.D(net288),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[10][5] ));
 DLH_X1 _10036_ (.D(net282),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[10][6] ));
 DLH_X1 _10037_ (.D(net276),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[10][7] ));
 DLH_X1 _10038_ (.D(net316),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[3][0] ));
 DLH_X1 _10039_ (.D(net313),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[3][1] ));
 DLH_X1 _10040_ (.D(net306),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[3][2] ));
 DLH_X1 _10041_ (.D(net298),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[3][3] ));
 DLH_X1 _10042_ (.D(net295),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[3][4] ));
 DLH_X1 _10043_ (.D(net288),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[3][5] ));
 DLH_X1 _10044_ (.D(net284),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[3][6] ));
 DLH_X1 _10045_ (.D(net276),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[3][7] ));
 DLH_X1 _10046_ (.D(net316),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[16][0] ));
 DLH_X1 _10047_ (.D(net312),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[16][1] ));
 DLH_X1 _10048_ (.D(net304),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[16][2] ));
 DLH_X1 _10049_ (.D(net298),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[16][3] ));
 DLH_X1 _10050_ (.D(net295),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[16][4] ));
 DLH_X1 _10051_ (.D(net292),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[16][5] ));
 DLH_X1 _10052_ (.D(net284),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[16][6] ));
 DLH_X1 _10053_ (.D(net276),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[16][7] ));
 DLH_X1 _10054_ (.D(net316),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[24][0] ));
 DLH_X1 _10055_ (.D(net313),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[24][1] ));
 DLH_X1 _10056_ (.D(net306),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[24][2] ));
 DLH_X1 _10057_ (.D(net298),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[24][3] ));
 DLH_X1 _10058_ (.D(net295),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[24][4] ));
 DLH_X1 _10059_ (.D(net292),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[24][5] ));
 DLH_X1 _10060_ (.D(net284),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[24][6] ));
 DLH_X1 _10061_ (.D(net277),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[24][7] ));
 DLH_X1 _10062_ (.D(net319),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[4][0] ));
 DLH_X1 _10063_ (.D(net313),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[4][1] ));
 DLH_X1 _10064_ (.D(net304),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[4][2] ));
 DLH_X1 _10065_ (.D(net298),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[4][3] ));
 DLH_X1 _10066_ (.D(net295),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[4][4] ));
 DLH_X1 _10067_ (.D(net292),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[4][5] ));
 DLH_X1 _10068_ (.D(net284),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[4][6] ));
 DLH_X1 _10069_ (.D(net276),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[4][7] ));
 DLH_X1 _10070_ (.D(net316),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[15][0] ));
 DLH_X1 _10071_ (.D(net313),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[15][1] ));
 DLH_X1 _10072_ (.D(net306),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[15][2] ));
 DLH_X1 _10073_ (.D(net303),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[15][3] ));
 DLH_X1 _10074_ (.D(net295),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[15][4] ));
 DLH_X1 _10075_ (.D(net288),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[15][5] ));
 DLH_X1 _10076_ (.D(net284),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[15][6] ));
 DLH_X1 _10077_ (.D(net276),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[15][7] ));
 DLH_X1 _10078_ (.D(net316),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[11][0] ));
 DLH_X1 _10079_ (.D(net313),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[11][1] ));
 DLH_X1 _10080_ (.D(net306),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[11][2] ));
 DLH_X1 _10081_ (.D(net298),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[11][3] ));
 DLH_X1 _10082_ (.D(net295),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[11][4] ));
 DLH_X1 _10083_ (.D(net288),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[11][5] ));
 DLH_X1 _10084_ (.D(net284),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[11][6] ));
 DLH_X1 _10085_ (.D(net277),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[11][7] ));
 DLH_X1 _10086_ (.D(net316),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[5][0] ));
 DLH_X1 _10087_ (.D(net313),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[5][1] ));
 DLH_X1 _10088_ (.D(net306),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[5][2] ));
 DLH_X1 _10089_ (.D(net298),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[5][3] ));
 DLH_X1 _10090_ (.D(net295),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[5][4] ));
 DLH_X1 _10091_ (.D(net288),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[5][5] ));
 DLH_X1 _10092_ (.D(net284),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[5][6] ));
 DLH_X1 _10093_ (.D(net276),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[5][7] ));
 DLH_X1 _10094_ (.D(net319),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[23][0] ));
 DLH_X1 _10095_ (.D(net313),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[23][1] ));
 DLH_X1 _10096_ (.D(net304),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[23][2] ));
 DLH_X1 _10097_ (.D(net298),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[23][3] ));
 DLH_X1 _10098_ (.D(net295),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[23][4] ));
 DLH_X1 _10099_ (.D(net288),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[23][5] ));
 DLH_X1 _10100_ (.D(net284),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[23][6] ));
 DLH_X1 _10101_ (.D(net276),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[23][7] ));
 DLH_X1 _10102_ (.D(net316),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[19][0] ));
 DLH_X1 _10103_ (.D(net313),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[19][1] ));
 DLH_X1 _10104_ (.D(net306),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[19][2] ));
 DLH_X1 _10105_ (.D(net298),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[19][3] ));
 DLH_X1 _10106_ (.D(net295),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[19][4] ));
 DLH_X1 _10107_ (.D(net288),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[19][5] ));
 DLH_X1 _10108_ (.D(net282),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[19][6] ));
 DLH_X1 _10109_ (.D(net277),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[19][7] ));
 DLH_X1 _10110_ (.D(net316),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[31][0] ));
 DLH_X1 _10111_ (.D(net313),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[31][1] ));
 DLH_X1 _10112_ (.D(net306),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[31][2] ));
 DLH_X1 _10113_ (.D(net298),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[31][3] ));
 DLH_X1 _10114_ (.D(net295),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[31][4] ));
 DLH_X1 _10115_ (.D(net288),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[31][5] ));
 DLH_X1 _10116_ (.D(net284),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[31][6] ));
 DLH_X1 _10117_ (.D(net276),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[31][7] ));
 DLH_X1 _10118_ (.D(net316),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[6][0] ));
 DLH_X1 _10119_ (.D(net313),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[6][1] ));
 DLH_X1 _10120_ (.D(net306),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[6][2] ));
 DLH_X1 _10121_ (.D(net303),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[6][3] ));
 DLH_X1 _10122_ (.D(net295),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[6][4] ));
 DLH_X1 _10123_ (.D(net288),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[6][5] ));
 DLH_X1 _10124_ (.D(net284),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[6][6] ));
 DLH_X1 _10125_ (.D(net276),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[6][7] ));
 DLH_X1 _10126_ (.D(net316),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[14][0] ));
 DLH_X1 _10127_ (.D(net312),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[14][1] ));
 DLH_X1 _10128_ (.D(net304),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[14][2] ));
 DLH_X1 _10129_ (.D(net298),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[14][3] ));
 DLH_X1 _10130_ (.D(net295),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[14][4] ));
 DLH_X1 _10131_ (.D(net292),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[14][5] ));
 DLH_X1 _10132_ (.D(net284),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[14][6] ));
 DLH_X1 _10133_ (.D(net279),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[14][7] ));
 DLH_X1 _10134_ (.D(net316),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[30][0] ));
 DLH_X1 _10135_ (.D(net313),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[30][1] ));
 DLH_X1 _10136_ (.D(net304),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[30][2] ));
 DLH_X1 _10137_ (.D(net298),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[30][3] ));
 DLH_X1 _10138_ (.D(net295),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[30][4] ));
 DLH_X1 _10139_ (.D(net292),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[30][5] ));
 DLH_X1 _10140_ (.D(net284),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[30][6] ));
 DLH_X1 _10141_ (.D(net279),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[30][7] ));
 DLH_X1 _10142_ (.D(net316),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[22][0] ));
 DLH_X1 _10143_ (.D(net313),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[22][1] ));
 DLH_X1 _10144_ (.D(net306),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[22][2] ));
 DLH_X1 _10145_ (.D(net298),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[22][3] ));
 DLH_X1 _10146_ (.D(net295),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[22][4] ));
 DLH_X1 _10147_ (.D(net292),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[22][5] ));
 DLH_X1 _10148_ (.D(net284),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[22][6] ));
 DLH_X1 _10149_ (.D(net276),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[22][7] ));
 DLH_X1 _10150_ (.D(net316),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[7][0] ));
 DLH_X1 _10151_ (.D(net313),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[7][1] ));
 DLH_X1 _10152_ (.D(net306),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[7][2] ));
 DLH_X1 _10153_ (.D(net298),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[7][3] ));
 DLH_X1 _10154_ (.D(net295),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[7][4] ));
 DLH_X1 _10155_ (.D(net288),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[7][5] ));
 DLH_X1 _10156_ (.D(net284),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[7][6] ));
 DLH_X1 _10157_ (.D(net276),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[7][7] ));
 DLH_X1 _10158_ (.D(net319),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[29][0] ));
 DLH_X1 _10159_ (.D(net313),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[29][1] ));
 DLH_X1 _10160_ (.D(net304),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[29][2] ));
 DLH_X1 _10161_ (.D(net298),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[29][3] ));
 DLH_X1 _10162_ (.D(net295),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[29][4] ));
 DLH_X1 _10163_ (.D(net292),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[29][5] ));
 DLH_X1 _10164_ (.D(net285),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[29][6] ));
 DLH_X1 _10165_ (.D(net279),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[29][7] ));
 DLH_X1 _10166_ (.D(net316),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[12][0] ));
 DLH_X1 _10167_ (.D(net313),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[12][1] ));
 DLH_X1 _10168_ (.D(net306),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[12][2] ));
 DLH_X1 _10169_ (.D(net303),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[12][3] ));
 DLH_X1 _10170_ (.D(net295),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[12][4] ));
 DLH_X1 _10171_ (.D(net288),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[12][5] ));
 DLH_X1 _10172_ (.D(net284),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[12][6] ));
 DLH_X1 _10173_ (.D(net277),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[12][7] ));
 DLH_X1 _10174_ (.D(net316),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[17][0] ));
 DLH_X1 _10175_ (.D(net313),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[17][1] ));
 DLH_X1 _10176_ (.D(net306),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[17][2] ));
 DLH_X1 _10177_ (.D(net303),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[17][3] ));
 DLH_X1 _10178_ (.D(net295),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[17][4] ));
 DLH_X1 _10179_ (.D(net288),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[17][5] ));
 DLH_X1 _10180_ (.D(net282),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[17][6] ));
 DLH_X1 _10181_ (.D(net276),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[17][7] ));
 DLH_X1 _10182_ (.D(net316),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[28][0] ));
 DLH_X1 _10183_ (.D(net313),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[28][1] ));
 DLH_X1 _10184_ (.D(net306),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[28][2] ));
 DLH_X1 _10185_ (.D(net303),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[28][3] ));
 DLH_X1 _10186_ (.D(net295),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[28][4] ));
 DLH_X1 _10187_ (.D(net288),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[28][5] ));
 DLH_X1 _10188_ (.D(net284),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[28][6] ));
 DLH_X1 _10189_ (.D(net276),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[28][7] ));
 DLH_X1 _10190_ (.D(net316),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[8][0] ));
 DLH_X1 _10191_ (.D(net313),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[8][1] ));
 DLH_X1 _10192_ (.D(net306),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[8][2] ));
 DLH_X1 _10193_ (.D(net298),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[8][3] ));
 DLH_X1 _10194_ (.D(net295),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[8][4] ));
 DLH_X1 _10195_ (.D(net288),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[8][5] ));
 DLH_X1 _10196_ (.D(net284),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[8][6] ));
 DLH_X1 _10197_ (.D(net277),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[8][7] ));
 DLH_X1 _10198_ (.D(net316),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[21][0] ));
 DLH_X1 _10199_ (.D(net313),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[21][1] ));
 DLH_X1 _10200_ (.D(net306),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[21][2] ));
 DLH_X1 _10201_ (.D(net298),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[21][3] ));
 DLH_X1 _10202_ (.D(net295),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[21][4] ));
 DLH_X1 _10203_ (.D(net288),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[21][5] ));
 DLH_X1 _10204_ (.D(net284),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[21][6] ));
 DLH_X1 _10205_ (.D(net276),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[21][7] ));
 DLH_X1 _10206_ (.D(net316),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[27][0] ));
 DLH_X1 _10207_ (.D(net313),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[27][1] ));
 DLH_X1 _10208_ (.D(net306),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[27][2] ));
 DLH_X1 _10209_ (.D(net303),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[27][3] ));
 DLH_X1 _10210_ (.D(net295),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[27][4] ));
 DLH_X1 _10211_ (.D(net288),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[27][5] ));
 DLH_X1 _10212_ (.D(net282),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[27][6] ));
 DLH_X1 _10213_ (.D(net277),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[27][7] ));
 DLH_X1 _10214_ (.D(net319),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[18][0] ));
 DLH_X1 _10215_ (.D(net313),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[18][1] ));
 DLH_X1 _10216_ (.D(net306),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[18][2] ));
 DLH_X1 _10217_ (.D(net303),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[18][3] ));
 DLH_X1 _10218_ (.D(net295),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[18][4] ));
 DLH_X1 _10219_ (.D(net288),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[18][5] ));
 DLH_X1 _10220_ (.D(net284),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[18][6] ));
 DLH_X1 _10221_ (.D(net277),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.mem[18][7] ));
 DLL_X1 _10222_ (.D(\lut.gen_sub_units_scm.__14.sub_unit_i.cg_we_global.en_i ),
    .GN(clknet_level_5_1_2116__00532_),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.cg_we_global.clk_en ));
 DLL_X1 _10223_ (.D(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__0.cg_i.en_i ),
    .GN(clknet_level_2_1_7137__00537_),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_en ));
 DLL_X1 _10224_ (.D(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__1.cg_i.en_i ),
    .GN(clknet_level_2_1_4128__00537_),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_en ));
 DLL_X1 _10225_ (.D(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__2.cg_i.en_i ),
    .GN(clknet_level_2_1_1119__00537_),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_en ));
 DLL_X1 _10226_ (.D(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__3.cg_i.en_i ),
    .GN(clknet_level_2_1_1119__00537_),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_en ));
 DLL_X1 _10227_ (.D(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__4.cg_i.en_i ),
    .GN(clknet_level_2_1_8140__00537_),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_en ));
 DLL_X1 _10228_ (.D(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__5.cg_i.en_i ),
    .GN(clknet_level_2_1_5131__00537_),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_en ));
 DLL_X1 _10229_ (.D(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__6.cg_i.en_i ),
    .GN(clknet_level_2_1_4128__00537_),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_en ));
 DLL_X1 _10230_ (.D(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__7.cg_i.en_i ),
    .GN(clknet_level_2_1_2122__00537_),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_en ));
 DLL_X1 _10231_ (.D(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__8.cg_i.en_i ),
    .GN(clknet_level_2_1_4128__00537_),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_en ));
 DLL_X1 _10232_ (.D(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__9.cg_i.en_i ),
    .GN(clknet_level_2_1_6134__00537_),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_en ));
 DLL_X1 _10233_ (.D(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__10.cg_i.en_i ),
    .GN(clknet_level_2_1_6134__00537_),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_en ));
 DLL_X1 _10234_ (.D(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__11.cg_i.en_i ),
    .GN(clknet_level_2_1_4128__00537_),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_en ));
 DLL_X1 _10235_ (.D(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__12.cg_i.en_i ),
    .GN(clknet_level_2_1_7137__00537_),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_en ));
 DLL_X1 _10236_ (.D(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__13.cg_i.en_i ),
    .GN(clknet_level_2_1_5131__00537_),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_en ));
 DLL_X1 _10237_ (.D(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__14.cg_i.en_i ),
    .GN(clknet_level_2_1_6134__00537_),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_en ));
 DLL_X1 _10238_ (.D(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__15.cg_i.en_i ),
    .GN(clknet_level_2_1_5131__00537_),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_en ));
 DLL_X1 _10239_ (.D(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__16.cg_i.en_i ),
    .GN(clknet_level_2_1_6134__00537_),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_en ));
 DLL_X1 _10240_ (.D(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__17.cg_i.en_i ),
    .GN(clknet_level_2_1_2122__00537_),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_en ));
 DLL_X1 _10241_ (.D(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__18.cg_i.en_i ),
    .GN(clknet_level_2_1_4128__00537_),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_en ));
 DLL_X1 _10242_ (.D(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__19.cg_i.en_i ),
    .GN(clknet_level_2_1_2122__00537_),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_en ));
 DLL_X1 _10243_ (.D(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__20.cg_i.en_i ),
    .GN(clknet_level_2_1_7137__00537_),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_en ));
 DLL_X1 _10244_ (.D(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__21.cg_i.en_i ),
    .GN(clknet_level_2_1_5131__00537_),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_en ));
 DLL_X1 _10245_ (.D(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__22.cg_i.en_i ),
    .GN(clknet_level_2_1_6134__00537_),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_en ));
 DLL_X1 _10246_ (.D(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__23.cg_i.en_i ),
    .GN(clknet_level_2_1_8140__00537_),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_en ));
 DLL_X1 _10247_ (.D(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__24.cg_i.en_i ),
    .GN(clknet_level_2_1_1119__00537_),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_en ));
 DLL_X1 _10248_ (.D(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__25.cg_i.en_i ),
    .GN(clknet_level_2_1_2122__00537_),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_en ));
 DLL_X1 _10249_ (.D(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__26.cg_i.en_i ),
    .GN(clknet_level_2_1_6134__00537_),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_en ));
 DLL_X1 _10250_ (.D(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__27.cg_i.en_i ),
    .GN(clknet_level_2_1_2122__00537_),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_en ));
 DLL_X1 _10251_ (.D(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__28.cg_i.en_i ),
    .GN(clknet_level_2_1_3125__00537_),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_en ));
 DLL_X1 _10252_ (.D(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__29.cg_i.en_i ),
    .GN(clknet_level_2_1_8140__00537_),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_en ));
 DLL_X1 _10253_ (.D(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__30.cg_i.en_i ),
    .GN(clknet_level_2_1_8140__00537_),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_en ));
 DLL_X1 _10254_ (.D(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__31.cg_i.en_i ),
    .GN(clknet_level_2_1_1119__00537_),
    .Q(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_en ));
 DLH_X1 _10255_ (.D(net320),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[13][0] ));
 DLH_X1 _10256_ (.D(net311),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[13][1] ));
 DLH_X1 _10257_ (.D(net305),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[13][2] ));
 DLH_X1 _10258_ (.D(net300),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[13][3] ));
 DLH_X1 _10259_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[4] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[13][4] ));
 DLH_X1 _10260_ (.D(net287),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[13][5] ));
 DLH_X1 _10261_ (.D(net285),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[13][6] ));
 DLH_X1 _10262_ (.D(net275),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[13][7] ));
 DLH_X1 _10263_ (.D(net317),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[1][0] ));
 DLH_X1 _10264_ (.D(net311),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[1][1] ));
 DLH_X1 _10265_ (.D(net306),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[1][2] ));
 DLH_X1 _10266_ (.D(net300),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[1][3] ));
 DLH_X1 _10267_ (.D(net294),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[1][4] ));
 DLH_X1 _10268_ (.D(net288),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[1][5] ));
 DLH_X1 _10269_ (.D(net285),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[1][6] ));
 DLH_X1 _10270_ (.D(net277),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[1][7] ));
 DLH_X1 _10271_ (.D(net320),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[26][0] ));
 DLH_X1 _10272_ (.D(net311),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[26][1] ));
 DLH_X1 _10273_ (.D(net305),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[26][2] ));
 DLH_X1 _10274_ (.D(net300),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[26][3] ));
 DLH_X1 _10275_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[4] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[26][4] ));
 DLH_X1 _10276_ (.D(net291),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[26][5] ));
 DLH_X1 _10277_ (.D(net285),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[26][6] ));
 DLH_X1 _10278_ (.D(net275),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[26][7] ));
 DLH_X1 _10279_ (.D(net320),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[9][0] ));
 DLH_X1 _10280_ (.D(net311),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[9][1] ));
 DLH_X1 _10281_ (.D(net305),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[9][2] ));
 DLH_X1 _10282_ (.D(net300),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[9][3] ));
 DLH_X1 _10283_ (.D(net294),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[9][4] ));
 DLH_X1 _10284_ (.D(net291),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[9][5] ));
 DLH_X1 _10285_ (.D(net283),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[9][6] ));
 DLH_X1 _10286_ (.D(net277),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[9][7] ));
 DLH_X1 _10287_ (.D(net317),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[0][0] ));
 DLH_X1 _10288_ (.D(net313),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[0][1] ));
 DLH_X1 _10289_ (.D(net306),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[0][2] ));
 DLH_X1 _10290_ (.D(net303),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[0][3] ));
 DLH_X1 _10291_ (.D(net294),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[0][4] ));
 DLH_X1 _10292_ (.D(net292),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[0][5] ));
 DLH_X1 _10293_ (.D(net285),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[0][6] ));
 DLH_X1 _10294_ (.D(net277),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[0][7] ));
 DLH_X1 _10295_ (.D(net317),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[20][0] ));
 DLH_X1 _10296_ (.D(net311),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[20][1] ));
 DLH_X1 _10297_ (.D(net305),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[20][2] ));
 DLH_X1 _10298_ (.D(net300),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[20][3] ));
 DLH_X1 _10299_ (.D(net294),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[20][4] ));
 DLH_X1 _10300_ (.D(net287),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[20][5] ));
 DLH_X1 _10301_ (.D(net285),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[20][6] ));
 DLH_X1 _10302_ (.D(net277),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[20][7] ));
 DLH_X1 _10303_ (.D(net317),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[2][0] ));
 DLH_X1 _10304_ (.D(net311),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[2][1] ));
 DLH_X1 _10305_ (.D(net305),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[2][2] ));
 DLH_X1 _10306_ (.D(net300),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[2][3] ));
 DLH_X1 _10307_ (.D(net294),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[2][4] ));
 DLH_X1 _10308_ (.D(net287),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[2][5] ));
 DLH_X1 _10309_ (.D(net285),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[2][6] ));
 DLH_X1 _10310_ (.D(net275),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[2][7] ));
 DLH_X1 _10311_ (.D(net317),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[25][0] ));
 DLH_X1 _10312_ (.D(net311),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[25][1] ));
 DLH_X1 _10313_ (.D(net305),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[25][2] ));
 DLH_X1 _10314_ (.D(net300),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[25][3] ));
 DLH_X1 _10315_ (.D(net294),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[25][4] ));
 DLH_X1 _10316_ (.D(net287),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[25][5] ));
 DLH_X1 _10317_ (.D(net285),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[25][6] ));
 DLH_X1 _10318_ (.D(net275),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[25][7] ));
 DLH_X1 _10319_ (.D(net317),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[10][0] ));
 DLH_X1 _10320_ (.D(net311),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[10][1] ));
 DLH_X1 _10321_ (.D(net306),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[10][2] ));
 DLH_X1 _10322_ (.D(net300),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[10][3] ));
 DLH_X1 _10323_ (.D(net294),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[10][4] ));
 DLH_X1 _10324_ (.D(net287),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[10][5] ));
 DLH_X1 _10325_ (.D(net285),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[10][6] ));
 DLH_X1 _10326_ (.D(net275),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[10][7] ));
 DLH_X1 _10327_ (.D(net317),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[3][0] ));
 DLH_X1 _10328_ (.D(net311),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[3][1] ));
 DLH_X1 _10329_ (.D(net306),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[3][2] ));
 DLH_X1 _10330_ (.D(net300),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[3][3] ));
 DLH_X1 _10331_ (.D(net294),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[3][4] ));
 DLH_X1 _10332_ (.D(net287),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[3][5] ));
 DLH_X1 _10333_ (.D(net285),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[3][6] ));
 DLH_X1 _10334_ (.D(net277),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[3][7] ));
 DLH_X1 _10335_ (.D(net317),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[16][0] ));
 DLH_X1 _10336_ (.D(net311),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[16][1] ));
 DLH_X1 _10337_ (.D(net305),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[16][2] ));
 DLH_X1 _10338_ (.D(net300),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[16][3] ));
 DLH_X1 _10339_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[4] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[16][4] ));
 DLH_X1 _10340_ (.D(net292),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[16][5] ));
 DLH_X1 _10341_ (.D(net285),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[16][6] ));
 DLH_X1 _10342_ (.D(net277),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[16][7] ));
 DLH_X1 _10343_ (.D(net317),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[24][0] ));
 DLH_X1 _10344_ (.D(net311),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[24][1] ));
 DLH_X1 _10345_ (.D(net305),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[24][2] ));
 DLH_X1 _10346_ (.D(net300),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[24][3] ));
 DLH_X1 _10347_ (.D(net294),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[24][4] ));
 DLH_X1 _10348_ (.D(net287),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[24][5] ));
 DLH_X1 _10349_ (.D(net284),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[24][6] ));
 DLH_X1 _10350_ (.D(net277),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[24][7] ));
 DLH_X1 _10351_ (.D(net320),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[4][0] ));
 DLH_X1 _10352_ (.D(net311),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[4][1] ));
 DLH_X1 _10353_ (.D(net305),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[4][2] ));
 DLH_X1 _10354_ (.D(net300),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[4][3] ));
 DLH_X1 _10355_ (.D(net294),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[4][4] ));
 DLH_X1 _10356_ (.D(net292),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[4][5] ));
 DLH_X1 _10357_ (.D(net284),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[4][6] ));
 DLH_X1 _10358_ (.D(net275),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[4][7] ));
 DLH_X1 _10359_ (.D(net317),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[15][0] ));
 DLH_X1 _10360_ (.D(net311),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[15][1] ));
 DLH_X1 _10361_ (.D(net306),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[15][2] ));
 DLH_X1 _10362_ (.D(net300),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[15][3] ));
 DLH_X1 _10363_ (.D(net294),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[15][4] ));
 DLH_X1 _10364_ (.D(net287),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[15][5] ));
 DLH_X1 _10365_ (.D(net284),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[15][6] ));
 DLH_X1 _10366_ (.D(net277),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[15][7] ));
 DLH_X1 _10367_ (.D(net320),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[11][0] ));
 DLH_X1 _10368_ (.D(net311),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[11][1] ));
 DLH_X1 _10369_ (.D(net306),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[11][2] ));
 DLH_X1 _10370_ (.D(net300),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[11][3] ));
 DLH_X1 _10371_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[4] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[11][4] ));
 DLH_X1 _10372_ (.D(net287),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[11][5] ));
 DLH_X1 _10373_ (.D(net284),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[11][6] ));
 DLH_X1 _10374_ (.D(net275),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[11][7] ));
 DLH_X1 _10375_ (.D(net317),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[5][0] ));
 DLH_X1 _10376_ (.D(net311),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[5][1] ));
 DLH_X1 _10377_ (.D(net305),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[5][2] ));
 DLH_X1 _10378_ (.D(net300),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[5][3] ));
 DLH_X1 _10379_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[4] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[5][4] ));
 DLH_X1 _10380_ (.D(net287),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[5][5] ));
 DLH_X1 _10381_ (.D(net285),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[5][6] ));
 DLH_X1 _10382_ (.D(net277),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[5][7] ));
 DLH_X1 _10383_ (.D(net317),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[23][0] ));
 DLH_X1 _10384_ (.D(net311),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[23][1] ));
 DLH_X1 _10385_ (.D(net305),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[23][2] ));
 DLH_X1 _10386_ (.D(net300),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[23][3] ));
 DLH_X1 _10387_ (.D(net294),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[23][4] ));
 DLH_X1 _10388_ (.D(net292),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[23][5] ));
 DLH_X1 _10389_ (.D(net285),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[23][6] ));
 DLH_X1 _10390_ (.D(net277),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[23][7] ));
 DLH_X1 _10391_ (.D(net317),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[19][0] ));
 DLH_X1 _10392_ (.D(net311),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[19][1] ));
 DLH_X1 _10393_ (.D(net306),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[19][2] ));
 DLH_X1 _10394_ (.D(net300),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[19][3] ));
 DLH_X1 _10395_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[4] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[19][4] ));
 DLH_X1 _10396_ (.D(net287),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[19][5] ));
 DLH_X1 _10397_ (.D(net285),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[19][6] ));
 DLH_X1 _10398_ (.D(net277),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[19][7] ));
 DLH_X1 _10399_ (.D(net317),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[31][0] ));
 DLH_X1 _10400_ (.D(net311),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[31][1] ));
 DLH_X1 _10401_ (.D(net306),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[31][2] ));
 DLH_X1 _10402_ (.D(net300),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[31][3] ));
 DLH_X1 _10403_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[4] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[31][4] ));
 DLH_X1 _10404_ (.D(net292),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[31][5] ));
 DLH_X1 _10405_ (.D(net284),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[31][6] ));
 DLH_X1 _10406_ (.D(net277),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[31][7] ));
 DLH_X1 _10407_ (.D(net317),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[6][0] ));
 DLH_X1 _10408_ (.D(net311),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[6][1] ));
 DLH_X1 _10409_ (.D(net305),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[6][2] ));
 DLH_X1 _10410_ (.D(net300),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[6][3] ));
 DLH_X1 _10411_ (.D(net294),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[6][4] ));
 DLH_X1 _10412_ (.D(net291),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[6][5] ));
 DLH_X1 _10413_ (.D(net285),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[6][6] ));
 DLH_X1 _10414_ (.D(net277),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[6][7] ));
 DLH_X1 _10415_ (.D(net317),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[14][0] ));
 DLH_X1 _10416_ (.D(net311),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[14][1] ));
 DLH_X1 _10417_ (.D(net306),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[14][2] ));
 DLH_X1 _10418_ (.D(net300),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[14][3] ));
 DLH_X1 _10419_ (.D(net294),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[14][4] ));
 DLH_X1 _10420_ (.D(net292),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[14][5] ));
 DLH_X1 _10421_ (.D(net284),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[14][6] ));
 DLH_X1 _10422_ (.D(net277),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[14][7] ));
 DLH_X1 _10423_ (.D(net317),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[30][0] ));
 DLH_X1 _10424_ (.D(net311),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[30][1] ));
 DLH_X1 _10425_ (.D(net306),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[30][2] ));
 DLH_X1 _10426_ (.D(net300),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[30][3] ));
 DLH_X1 _10427_ (.D(net294),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[30][4] ));
 DLH_X1 _10428_ (.D(net287),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[30][5] ));
 DLH_X1 _10429_ (.D(net284),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[30][6] ));
 DLH_X1 _10430_ (.D(net277),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[30][7] ));
 DLH_X1 _10431_ (.D(net317),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[22][0] ));
 DLH_X1 _10432_ (.D(net311),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[22][1] ));
 DLH_X1 _10433_ (.D(net305),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[22][2] ));
 DLH_X1 _10434_ (.D(net300),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[22][3] ));
 DLH_X1 _10435_ (.D(net294),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[22][4] ));
 DLH_X1 _10436_ (.D(net287),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[22][5] ));
 DLH_X1 _10437_ (.D(net285),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[22][6] ));
 DLH_X1 _10438_ (.D(net275),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[22][7] ));
 DLH_X1 _10439_ (.D(net317),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[7][0] ));
 DLH_X1 _10440_ (.D(net311),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[7][1] ));
 DLH_X1 _10441_ (.D(net305),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[7][2] ));
 DLH_X1 _10442_ (.D(net300),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[7][3] ));
 DLH_X1 _10443_ (.D(net294),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[7][4] ));
 DLH_X1 _10444_ (.D(net287),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[7][5] ));
 DLH_X1 _10445_ (.D(net285),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[7][6] ));
 DLH_X1 _10446_ (.D(net277),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[7][7] ));
 DLH_X1 _10447_ (.D(net320),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[29][0] ));
 DLH_X1 _10448_ (.D(net311),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[29][1] ));
 DLH_X1 _10449_ (.D(net306),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[29][2] ));
 DLH_X1 _10450_ (.D(net300),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[29][3] ));
 DLH_X1 _10451_ (.D(net294),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[29][4] ));
 DLH_X1 _10452_ (.D(net292),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[29][5] ));
 DLH_X1 _10453_ (.D(net285),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[29][6] ));
 DLH_X1 _10454_ (.D(net277),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[29][7] ));
 DLH_X1 _10455_ (.D(net317),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[12][0] ));
 DLH_X1 _10456_ (.D(net311),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[12][1] ));
 DLH_X1 _10457_ (.D(net305),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[12][2] ));
 DLH_X1 _10458_ (.D(net300),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[12][3] ));
 DLH_X1 _10459_ (.D(net294),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[12][4] ));
 DLH_X1 _10460_ (.D(net292),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[12][5] ));
 DLH_X1 _10461_ (.D(net285),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[12][6] ));
 DLH_X1 _10462_ (.D(net277),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[12][7] ));
 DLH_X1 _10463_ (.D(net317),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[17][0] ));
 DLH_X1 _10464_ (.D(net311),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[17][1] ));
 DLH_X1 _10465_ (.D(net306),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[17][2] ));
 DLH_X1 _10466_ (.D(net300),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[17][3] ));
 DLH_X1 _10467_ (.D(net294),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[17][4] ));
 DLH_X1 _10468_ (.D(net287),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[17][5] ));
 DLH_X1 _10469_ (.D(net285),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[17][6] ));
 DLH_X1 _10470_ (.D(net277),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[17][7] ));
 DLH_X1 _10471_ (.D(net317),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[28][0] ));
 DLH_X1 _10472_ (.D(net311),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[28][1] ));
 DLH_X1 _10473_ (.D(net306),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[28][2] ));
 DLH_X1 _10474_ (.D(net300),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[28][3] ));
 DLH_X1 _10475_ (.D(net294),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[28][4] ));
 DLH_X1 _10476_ (.D(net292),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[28][5] ));
 DLH_X1 _10477_ (.D(net284),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[28][6] ));
 DLH_X1 _10478_ (.D(net277),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[28][7] ));
 DLH_X1 _10479_ (.D(net320),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[8][0] ));
 DLH_X1 _10480_ (.D(net311),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[8][1] ));
 DLH_X1 _10481_ (.D(net306),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[8][2] ));
 DLH_X1 _10482_ (.D(net300),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[8][3] ));
 DLH_X1 _10483_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[4] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[8][4] ));
 DLH_X1 _10484_ (.D(net291),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[8][5] ));
 DLH_X1 _10485_ (.D(net285),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[8][6] ));
 DLH_X1 _10486_ (.D(net277),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[8][7] ));
 DLH_X1 _10487_ (.D(net317),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[21][0] ));
 DLH_X1 _10488_ (.D(net311),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[21][1] ));
 DLH_X1 _10489_ (.D(net305),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[21][2] ));
 DLH_X1 _10490_ (.D(net300),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[21][3] ));
 DLH_X1 _10491_ (.D(net294),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[21][4] ));
 DLH_X1 _10492_ (.D(net292),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[21][5] ));
 DLH_X1 _10493_ (.D(net284),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[21][6] ));
 DLH_X1 _10494_ (.D(net277),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[21][7] ));
 DLH_X1 _10495_ (.D(net317),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[27][0] ));
 DLH_X1 _10496_ (.D(net311),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[27][1] ));
 DLH_X1 _10497_ (.D(net306),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[27][2] ));
 DLH_X1 _10498_ (.D(net300),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[27][3] ));
 DLH_X1 _10499_ (.D(net294),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[27][4] ));
 DLH_X1 _10500_ (.D(net287),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[27][5] ));
 DLH_X1 _10501_ (.D(net284),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[27][6] ));
 DLH_X1 _10502_ (.D(net277),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[27][7] ));
 DLH_X1 _10503_ (.D(net320),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[18][0] ));
 DLH_X1 _10504_ (.D(net311),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[18][1] ));
 DLH_X1 _10505_ (.D(net305),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[18][2] ));
 DLH_X1 _10506_ (.D(net300),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[18][3] ));
 DLH_X1 _10507_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[4] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[18][4] ));
 DLH_X1 _10508_ (.D(net287),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[18][5] ));
 DLH_X1 _10509_ (.D(net285),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[18][6] ));
 DLH_X1 _10510_ (.D(net277),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.mem[18][7] ));
 DLL_X1 _10511_ (.D(\lut.gen_sub_units_scm.__13.sub_unit_i.cg_we_global.en_i ),
    .GN(clknet_level_5_1_4320__00532_),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.cg_we_global.clk_en ));
 DLL_X1 _10512_ (.D(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__0.cg_i.en_i ),
    .GN(clknet_level_2_1_5335__00540_),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_en ));
 DLL_X1 _10513_ (.D(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__1.cg_i.en_i ),
    .GN(clknet_level_2_1_8344__00540_),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_en ));
 DLL_X1 _10514_ (.D(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__2.cg_i.en_i ),
    .GN(clknet_level_2_1_3329__00540_),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_en ));
 DLL_X1 _10515_ (.D(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__3.cg_i.en_i ),
    .GN(clknet_level_2_1_6338__00540_),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_en ));
 DLL_X1 _10516_ (.D(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__4.cg_i.en_i ),
    .GN(clknet_level_2_1_4332__00540_),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_en ));
 DLL_X1 _10517_ (.D(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__5.cg_i.en_i ),
    .GN(clknet_level_2_1_3329__00540_),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_en ));
 DLL_X1 _10518_ (.D(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__6.cg_i.en_i ),
    .GN(clknet_level_2_1_3329__00540_),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_en ));
 DLL_X1 _10519_ (.D(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__7.cg_i.en_i ),
    .GN(clknet_level_2_1_1323__00540_),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_en ));
 DLL_X1 _10520_ (.D(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__8.cg_i.en_i ),
    .GN(clknet_level_2_1_7341__00540_),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_en ));
 DLL_X1 _10521_ (.D(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__9.cg_i.en_i ),
    .GN(clknet_level_2_1_4332__00540_),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_en ));
 DLL_X1 _10522_ (.D(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__10.cg_i.en_i ),
    .GN(clknet_level_2_1_8344__00540_),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_en ));
 DLL_X1 _10523_ (.D(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__11.cg_i.en_i ),
    .GN(clknet_level_2_1_4332__00540_),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_en ));
 DLL_X1 _10524_ (.D(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__12.cg_i.en_i ),
    .GN(clknet_level_2_1_2326__00540_),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_en ));
 DLL_X1 _10525_ (.D(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__13.cg_i.en_i ),
    .GN(clknet_level_2_1_3329__00540_),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_en ));
 DLL_X1 _10526_ (.D(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__14.cg_i.en_i ),
    .GN(clknet_level_2_1_5335__00540_),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_en ));
 DLL_X1 _10527_ (.D(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__15.cg_i.en_i ),
    .GN(clknet_level_2_1_1323__00540_),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_en ));
 DLL_X1 _10528_ (.D(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__16.cg_i.en_i ),
    .GN(clknet_level_2_1_8344__00540_),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_en ));
 DLL_X1 _10529_ (.D(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__17.cg_i.en_i ),
    .GN(clknet_level_2_1_5335__00540_),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_en ));
 DLL_X1 _10530_ (.D(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__18.cg_i.en_i ),
    .GN(clknet_level_2_1_7341__00540_),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_en ));
 DLL_X1 _10531_ (.D(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__19.cg_i.en_i ),
    .GN(clknet_level_2_1_4332__00540_),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_en ));
 DLL_X1 _10532_ (.D(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__20.cg_i.en_i ),
    .GN(clknet_level_2_1_1323__00540_),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_en ));
 DLL_X1 _10533_ (.D(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__21.cg_i.en_i ),
    .GN(clknet_level_2_1_1323__00540_),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_en ));
 DLL_X1 _10534_ (.D(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__22.cg_i.en_i ),
    .GN(clknet_level_2_1_4332__00540_),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_en ));
 DLL_X1 _10535_ (.D(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__23.cg_i.en_i ),
    .GN(clknet_level_2_1_7341__00540_),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_en ));
 DLL_X1 _10536_ (.D(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__24.cg_i.en_i ),
    .GN(clknet_level_2_1_3329__00540_),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_en ));
 DLL_X1 _10537_ (.D(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__25.cg_i.en_i ),
    .GN(clknet_level_2_1_1323__00540_),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_en ));
 DLL_X1 _10538_ (.D(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__26.cg_i.en_i ),
    .GN(clknet_level_2_1_3329__00540_),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_en ));
 DLL_X1 _10539_ (.D(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__27.cg_i.en_i ),
    .GN(clknet_level_2_1_2326__00540_),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_en ));
 DLL_X1 _10540_ (.D(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__28.cg_i.en_i ),
    .GN(clknet_level_2_1_6338__00540_),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_en ));
 DLL_X1 _10541_ (.D(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__29.cg_i.en_i ),
    .GN(clknet_level_2_1_8344__00540_),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_en ));
 DLL_X1 _10542_ (.D(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__30.cg_i.en_i ),
    .GN(clknet_level_2_1_2326__00540_),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_en ));
 DLL_X1 _10543_ (.D(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__31.cg_i.en_i ),
    .GN(clknet_level_2_1_6338__00540_),
    .Q(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_en ));
 DLH_X1 _10544_ (.D(net318),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[13][0] ));
 DLH_X1 _10545_ (.D(net314),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[13][1] ));
 DLH_X1 _10546_ (.D(net309),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[13][2] ));
 DLH_X1 _10547_ (.D(net301),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[13][3] ));
 DLH_X1 _10548_ (.D(net296),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[13][4] ));
 DLH_X1 _10549_ (.D(net289),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[13][5] ));
 DLH_X1 _10550_ (.D(net281),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[13][6] ));
 DLH_X1 _10551_ (.D(net278),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[13][7] ));
 DLH_X1 _10552_ (.D(net318),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[1][0] ));
 DLH_X1 _10553_ (.D(net314),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[1][1] ));
 DLH_X1 _10554_ (.D(net309),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[1][2] ));
 DLH_X1 _10555_ (.D(net301),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[1][3] ));
 DLH_X1 _10556_ (.D(net296),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[1][4] ));
 DLH_X1 _10557_ (.D(net289),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[1][5] ));
 DLH_X1 _10558_ (.D(net281),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[1][6] ));
 DLH_X1 _10559_ (.D(net278),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[1][7] ));
 DLH_X1 _10560_ (.D(net318),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[26][0] ));
 DLH_X1 _10561_ (.D(net314),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[26][1] ));
 DLH_X1 _10562_ (.D(net309),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[26][2] ));
 DLH_X1 _10563_ (.D(net301),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[26][3] ));
 DLH_X1 _10564_ (.D(net296),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[26][4] ));
 DLH_X1 _10565_ (.D(net289),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[26][5] ));
 DLH_X1 _10566_ (.D(net281),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[26][6] ));
 DLH_X1 _10567_ (.D(net278),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[26][7] ));
 DLH_X1 _10568_ (.D(net318),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[9][0] ));
 DLH_X1 _10569_ (.D(net314),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[9][1] ));
 DLH_X1 _10570_ (.D(net309),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[9][2] ));
 DLH_X1 _10571_ (.D(net301),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[9][3] ));
 DLH_X1 _10572_ (.D(net296),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[9][4] ));
 DLH_X1 _10573_ (.D(net289),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[9][5] ));
 DLH_X1 _10574_ (.D(net281),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[9][6] ));
 DLH_X1 _10575_ (.D(net278),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[9][7] ));
 DLH_X1 _10576_ (.D(net319),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[0][0] ));
 DLH_X1 _10577_ (.D(net313),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[0][1] ));
 DLH_X1 _10578_ (.D(net304),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[0][2] ));
 DLH_X1 _10579_ (.D(net303),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[0][3] ));
 DLH_X1 _10580_ (.D(net295),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[0][4] ));
 DLH_X1 _10581_ (.D(net292),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[0][5] ));
 DLH_X1 _10582_ (.D(net281),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[0][6] ));
 DLH_X1 _10583_ (.D(net279),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[0][7] ));
 DLH_X1 _10584_ (.D(net318),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[20][0] ));
 DLH_X1 _10585_ (.D(net314),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[20][1] ));
 DLH_X1 _10586_ (.D(net309),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[20][2] ));
 DLH_X1 _10587_ (.D(net301),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[20][3] ));
 DLH_X1 _10588_ (.D(net296),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[20][4] ));
 DLH_X1 _10589_ (.D(net289),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[20][5] ));
 DLH_X1 _10590_ (.D(net281),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[20][6] ));
 DLH_X1 _10591_ (.D(net278),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[20][7] ));
 DLH_X1 _10592_ (.D(net318),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[2][0] ));
 DLH_X1 _10593_ (.D(net314),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[2][1] ));
 DLH_X1 _10594_ (.D(net309),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[2][2] ));
 DLH_X1 _10595_ (.D(net301),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[2][3] ));
 DLH_X1 _10596_ (.D(net296),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[2][4] ));
 DLH_X1 _10597_ (.D(net289),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[2][5] ));
 DLH_X1 _10598_ (.D(net281),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[2][6] ));
 DLH_X1 _10599_ (.D(net278),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[2][7] ));
 DLH_X1 _10600_ (.D(net318),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[25][0] ));
 DLH_X1 _10601_ (.D(net314),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[25][1] ));
 DLH_X1 _10602_ (.D(net309),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[25][2] ));
 DLH_X1 _10603_ (.D(net301),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[25][3] ));
 DLH_X1 _10604_ (.D(net296),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[25][4] ));
 DLH_X1 _10605_ (.D(net289),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[25][5] ));
 DLH_X1 _10606_ (.D(net281),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[25][6] ));
 DLH_X1 _10607_ (.D(net278),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[25][7] ));
 DLH_X1 _10608_ (.D(net318),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[10][0] ));
 DLH_X1 _10609_ (.D(net314),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[10][1] ));
 DLH_X1 _10610_ (.D(net309),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[10][2] ));
 DLH_X1 _10611_ (.D(net301),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[10][3] ));
 DLH_X1 _10612_ (.D(net296),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[10][4] ));
 DLH_X1 _10613_ (.D(net289),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[10][5] ));
 DLH_X1 _10614_ (.D(net281),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[10][6] ));
 DLH_X1 _10615_ (.D(net278),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[10][7] ));
 DLH_X1 _10616_ (.D(net318),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[3][0] ));
 DLH_X1 _10617_ (.D(net314),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[3][1] ));
 DLH_X1 _10618_ (.D(net309),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[3][2] ));
 DLH_X1 _10619_ (.D(net301),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[3][3] ));
 DLH_X1 _10620_ (.D(net296),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[3][4] ));
 DLH_X1 _10621_ (.D(net289),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[3][5] ));
 DLH_X1 _10622_ (.D(net281),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[3][6] ));
 DLH_X1 _10623_ (.D(net278),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[3][7] ));
 DLH_X1 _10624_ (.D(net318),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[16][0] ));
 DLH_X1 _10625_ (.D(net314),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[16][1] ));
 DLH_X1 _10626_ (.D(net309),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[16][2] ));
 DLH_X1 _10627_ (.D(net301),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[16][3] ));
 DLH_X1 _10628_ (.D(net296),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[16][4] ));
 DLH_X1 _10629_ (.D(net289),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[16][5] ));
 DLH_X1 _10630_ (.D(net281),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[16][6] ));
 DLH_X1 _10631_ (.D(net278),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[16][7] ));
 DLH_X1 _10632_ (.D(net318),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[24][0] ));
 DLH_X1 _10633_ (.D(net314),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[24][1] ));
 DLH_X1 _10634_ (.D(net309),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[24][2] ));
 DLH_X1 _10635_ (.D(net301),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[24][3] ));
 DLH_X1 _10636_ (.D(net296),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[24][4] ));
 DLH_X1 _10637_ (.D(net289),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[24][5] ));
 DLH_X1 _10638_ (.D(net281),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[24][6] ));
 DLH_X1 _10639_ (.D(net278),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[24][7] ));
 DLH_X1 _10640_ (.D(net318),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[4][0] ));
 DLH_X1 _10641_ (.D(net314),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[4][1] ));
 DLH_X1 _10642_ (.D(net309),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[4][2] ));
 DLH_X1 _10643_ (.D(net301),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[4][3] ));
 DLH_X1 _10644_ (.D(net296),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[4][4] ));
 DLH_X1 _10645_ (.D(net289),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[4][5] ));
 DLH_X1 _10646_ (.D(net281),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[4][6] ));
 DLH_X1 _10647_ (.D(net278),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[4][7] ));
 DLH_X1 _10648_ (.D(net318),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[15][0] ));
 DLH_X1 _10649_ (.D(net314),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[15][1] ));
 DLH_X1 _10650_ (.D(net309),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[15][2] ));
 DLH_X1 _10651_ (.D(net301),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[15][3] ));
 DLH_X1 _10652_ (.D(net296),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[15][4] ));
 DLH_X1 _10653_ (.D(net289),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[15][5] ));
 DLH_X1 _10654_ (.D(net281),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[15][6] ));
 DLH_X1 _10655_ (.D(net278),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[15][7] ));
 DLH_X1 _10656_ (.D(net318),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[11][0] ));
 DLH_X1 _10657_ (.D(net314),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[11][1] ));
 DLH_X1 _10658_ (.D(net309),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[11][2] ));
 DLH_X1 _10659_ (.D(net301),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[11][3] ));
 DLH_X1 _10660_ (.D(net296),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[11][4] ));
 DLH_X1 _10661_ (.D(net289),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[11][5] ));
 DLH_X1 _10662_ (.D(net281),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[11][6] ));
 DLH_X1 _10663_ (.D(net278),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[11][7] ));
 DLH_X1 _10664_ (.D(net318),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[5][0] ));
 DLH_X1 _10665_ (.D(net314),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[5][1] ));
 DLH_X1 _10666_ (.D(net309),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[5][2] ));
 DLH_X1 _10667_ (.D(net301),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[5][3] ));
 DLH_X1 _10668_ (.D(net296),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[5][4] ));
 DLH_X1 _10669_ (.D(net289),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[5][5] ));
 DLH_X1 _10670_ (.D(net281),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[5][6] ));
 DLH_X1 _10671_ (.D(net278),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[5][7] ));
 DLH_X1 _10672_ (.D(net318),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[23][0] ));
 DLH_X1 _10673_ (.D(net314),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[23][1] ));
 DLH_X1 _10674_ (.D(net309),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[23][2] ));
 DLH_X1 _10675_ (.D(net301),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[23][3] ));
 DLH_X1 _10676_ (.D(net296),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[23][4] ));
 DLH_X1 _10677_ (.D(net289),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[23][5] ));
 DLH_X1 _10678_ (.D(net281),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[23][6] ));
 DLH_X1 _10679_ (.D(net278),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[23][7] ));
 DLH_X1 _10680_ (.D(net318),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[19][0] ));
 DLH_X1 _10681_ (.D(net314),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[19][1] ));
 DLH_X1 _10682_ (.D(net309),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[19][2] ));
 DLH_X1 _10683_ (.D(net301),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[19][3] ));
 DLH_X1 _10684_ (.D(net296),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[19][4] ));
 DLH_X1 _10685_ (.D(net289),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[19][5] ));
 DLH_X1 _10686_ (.D(net281),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[19][6] ));
 DLH_X1 _10687_ (.D(net278),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[19][7] ));
 DLH_X1 _10688_ (.D(net318),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[31][0] ));
 DLH_X1 _10689_ (.D(net314),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[31][1] ));
 DLH_X1 _10690_ (.D(net309),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[31][2] ));
 DLH_X1 _10691_ (.D(net301),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[31][3] ));
 DLH_X1 _10692_ (.D(net296),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[31][4] ));
 DLH_X1 _10693_ (.D(net289),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[31][5] ));
 DLH_X1 _10694_ (.D(net281),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[31][6] ));
 DLH_X1 _10695_ (.D(net278),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[31][7] ));
 DLH_X1 _10696_ (.D(net318),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[6][0] ));
 DLH_X1 _10697_ (.D(net314),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[6][1] ));
 DLH_X1 _10698_ (.D(net309),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[6][2] ));
 DLH_X1 _10699_ (.D(net301),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[6][3] ));
 DLH_X1 _10700_ (.D(net296),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[6][4] ));
 DLH_X1 _10701_ (.D(net289),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[6][5] ));
 DLH_X1 _10702_ (.D(net281),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[6][6] ));
 DLH_X1 _10703_ (.D(net278),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[6][7] ));
 DLH_X1 _10704_ (.D(net318),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[14][0] ));
 DLH_X1 _10705_ (.D(net314),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[14][1] ));
 DLH_X1 _10706_ (.D(net309),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[14][2] ));
 DLH_X1 _10707_ (.D(net301),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[14][3] ));
 DLH_X1 _10708_ (.D(net296),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[14][4] ));
 DLH_X1 _10709_ (.D(net289),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[14][5] ));
 DLH_X1 _10710_ (.D(net281),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[14][6] ));
 DLH_X1 _10711_ (.D(net278),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[14][7] ));
 DLH_X1 _10712_ (.D(net318),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[30][0] ));
 DLH_X1 _10713_ (.D(net314),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[30][1] ));
 DLH_X1 _10714_ (.D(net309),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[30][2] ));
 DLH_X1 _10715_ (.D(net301),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[30][3] ));
 DLH_X1 _10716_ (.D(net296),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[30][4] ));
 DLH_X1 _10717_ (.D(net289),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[30][5] ));
 DLH_X1 _10718_ (.D(net281),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[30][6] ));
 DLH_X1 _10719_ (.D(net278),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[30][7] ));
 DLH_X1 _10720_ (.D(net318),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[22][0] ));
 DLH_X1 _10721_ (.D(net314),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[22][1] ));
 DLH_X1 _10722_ (.D(net309),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[22][2] ));
 DLH_X1 _10723_ (.D(net301),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[22][3] ));
 DLH_X1 _10724_ (.D(net296),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[22][4] ));
 DLH_X1 _10725_ (.D(net289),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[22][5] ));
 DLH_X1 _10726_ (.D(net281),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[22][6] ));
 DLH_X1 _10727_ (.D(net278),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[22][7] ));
 DLH_X1 _10728_ (.D(net318),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[7][0] ));
 DLH_X1 _10729_ (.D(net314),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[7][1] ));
 DLH_X1 _10730_ (.D(net309),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[7][2] ));
 DLH_X1 _10731_ (.D(net301),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[7][3] ));
 DLH_X1 _10732_ (.D(net296),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[7][4] ));
 DLH_X1 _10733_ (.D(net289),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[7][5] ));
 DLH_X1 _10734_ (.D(net281),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[7][6] ));
 DLH_X1 _10735_ (.D(net278),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[7][7] ));
 DLH_X1 _10736_ (.D(net318),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[29][0] ));
 DLH_X1 _10737_ (.D(net314),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[29][1] ));
 DLH_X1 _10738_ (.D(net309),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[29][2] ));
 DLH_X1 _10739_ (.D(net301),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[29][3] ));
 DLH_X1 _10740_ (.D(net296),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[29][4] ));
 DLH_X1 _10741_ (.D(net289),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[29][5] ));
 DLH_X1 _10742_ (.D(net281),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[29][6] ));
 DLH_X1 _10743_ (.D(net278),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[29][7] ));
 DLH_X1 _10744_ (.D(net318),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[12][0] ));
 DLH_X1 _10745_ (.D(net314),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[12][1] ));
 DLH_X1 _10746_ (.D(net309),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[12][2] ));
 DLH_X1 _10747_ (.D(net301),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[12][3] ));
 DLH_X1 _10748_ (.D(net296),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[12][4] ));
 DLH_X1 _10749_ (.D(net289),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[12][5] ));
 DLH_X1 _10750_ (.D(net281),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[12][6] ));
 DLH_X1 _10751_ (.D(net278),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[12][7] ));
 DLH_X1 _10752_ (.D(net318),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[17][0] ));
 DLH_X1 _10753_ (.D(net314),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[17][1] ));
 DLH_X1 _10754_ (.D(net309),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[17][2] ));
 DLH_X1 _10755_ (.D(net301),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[17][3] ));
 DLH_X1 _10756_ (.D(net296),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[17][4] ));
 DLH_X1 _10757_ (.D(net289),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[17][5] ));
 DLH_X1 _10758_ (.D(net281),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[17][6] ));
 DLH_X1 _10759_ (.D(net278),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[17][7] ));
 DLH_X1 _10760_ (.D(net318),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[28][0] ));
 DLH_X1 _10761_ (.D(net314),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[28][1] ));
 DLH_X1 _10762_ (.D(net309),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[28][2] ));
 DLH_X1 _10763_ (.D(net301),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[28][3] ));
 DLH_X1 _10764_ (.D(net296),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[28][4] ));
 DLH_X1 _10765_ (.D(net289),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[28][5] ));
 DLH_X1 _10766_ (.D(net281),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[28][6] ));
 DLH_X1 _10767_ (.D(net278),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[28][7] ));
 DLH_X1 _10768_ (.D(net318),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[8][0] ));
 DLH_X1 _10769_ (.D(net314),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[8][1] ));
 DLH_X1 _10770_ (.D(net309),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[8][2] ));
 DLH_X1 _10771_ (.D(net301),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[8][3] ));
 DLH_X1 _10772_ (.D(net296),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[8][4] ));
 DLH_X1 _10773_ (.D(net289),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[8][5] ));
 DLH_X1 _10774_ (.D(net281),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[8][6] ));
 DLH_X1 _10775_ (.D(net278),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[8][7] ));
 DLH_X1 _10776_ (.D(net318),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[21][0] ));
 DLH_X1 _10777_ (.D(net314),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[21][1] ));
 DLH_X1 _10778_ (.D(net309),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[21][2] ));
 DLH_X1 _10779_ (.D(net301),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[21][3] ));
 DLH_X1 _10780_ (.D(net296),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[21][4] ));
 DLH_X1 _10781_ (.D(net289),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[21][5] ));
 DLH_X1 _10782_ (.D(net281),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[21][6] ));
 DLH_X1 _10783_ (.D(net278),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[21][7] ));
 DLH_X1 _10784_ (.D(net318),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[27][0] ));
 DLH_X1 _10785_ (.D(net314),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[27][1] ));
 DLH_X1 _10786_ (.D(net309),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[27][2] ));
 DLH_X1 _10787_ (.D(net301),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[27][3] ));
 DLH_X1 _10788_ (.D(net296),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[27][4] ));
 DLH_X1 _10789_ (.D(net289),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[27][5] ));
 DLH_X1 _10790_ (.D(net281),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[27][6] ));
 DLH_X1 _10791_ (.D(net278),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[27][7] ));
 DLH_X1 _10792_ (.D(net318),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[18][0] ));
 DLH_X1 _10793_ (.D(net314),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[18][1] ));
 DLH_X1 _10794_ (.D(net309),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[18][2] ));
 DLH_X1 _10795_ (.D(net301),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[18][3] ));
 DLH_X1 _10796_ (.D(net296),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[18][4] ));
 DLH_X1 _10797_ (.D(net289),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[18][5] ));
 DLH_X1 _10798_ (.D(net281),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[18][6] ));
 DLH_X1 _10799_ (.D(net278),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.mem[18][7] ));
 DLL_X1 _10800_ (.D(\lut.gen_sub_units_scm.__12.sub_unit_i.cg_we_global.en_i ),
    .GN(clknet_level_5_1_2116__00532_),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.cg_we_global.clk_en ));
 DLL_X1 _10801_ (.D(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__0.cg_i.en_i ),
    .GN(clknet_level_2_1_6158__00543_),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_en ));
 DLL_X1 _10802_ (.D(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__1.cg_i.en_i ),
    .GN(clknet_level_2_1_8164__00543_),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_en ));
 DLL_X1 _10803_ (.D(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__2.cg_i.en_i ),
    .GN(clknet_level_2_1_6158__00543_),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_en ));
 DLL_X1 _10804_ (.D(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__3.cg_i.en_i ),
    .GN(clknet_level_2_1_8164__00543_),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_en ));
 DLL_X1 _10805_ (.D(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__4.cg_i.en_i ),
    .GN(clknet_level_2_1_3149__00543_),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_en ));
 DLL_X1 _10806_ (.D(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__5.cg_i.en_i ),
    .GN(clknet_level_2_1_1143__00543_),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_en ));
 DLL_X1 _10807_ (.D(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__6.cg_i.en_i ),
    .GN(clknet_level_2_1_4152__00543_),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_en ));
 DLL_X1 _10808_ (.D(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__7.cg_i.en_i ),
    .GN(clknet_level_2_1_4152__00543_),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_en ));
 DLL_X1 _10809_ (.D(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__8.cg_i.en_i ),
    .GN(clknet_level_2_1_3149__00543_),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_en ));
 DLL_X1 _10810_ (.D(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__9.cg_i.en_i ),
    .GN(clknet_level_2_1_4152__00543_),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_en ));
 DLL_X1 _10811_ (.D(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__10.cg_i.en_i ),
    .GN(clknet_level_2_1_7161__00543_),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_en ));
 DLL_X1 _10812_ (.D(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__11.cg_i.en_i ),
    .GN(clknet_level_2_1_4152__00543_),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_en ));
 DLL_X1 _10813_ (.D(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__12.cg_i.en_i ),
    .GN(clknet_level_2_1_5155__00543_),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_en ));
 DLL_X1 _10814_ (.D(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__13.cg_i.en_i ),
    .GN(clknet_level_2_1_3149__00543_),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_en ));
 DLL_X1 _10815_ (.D(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__14.cg_i.en_i ),
    .GN(clknet_level_2_1_6158__00543_),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_en ));
 DLL_X1 _10816_ (.D(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__15.cg_i.en_i ),
    .GN(clknet_level_2_1_4152__00543_),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_en ));
 DLL_X1 _10817_ (.D(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__16.cg_i.en_i ),
    .GN(clknet_level_2_1_8164__00543_),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_en ));
 DLL_X1 _10818_ (.D(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__17.cg_i.en_i ),
    .GN(clknet_level_2_1_5155__00543_),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_en ));
 DLL_X1 _10819_ (.D(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__18.cg_i.en_i ),
    .GN(clknet_level_2_1_2146__00543_),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_en ));
 DLL_X1 _10820_ (.D(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__19.cg_i.en_i ),
    .GN(clknet_level_2_1_7161__00543_),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_en ));
 DLL_X1 _10821_ (.D(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__20.cg_i.en_i ),
    .GN(clknet_level_2_1_7161__00543_),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_en ));
 DLL_X1 _10822_ (.D(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__21.cg_i.en_i ),
    .GN(clknet_level_2_1_4152__00543_),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_en ));
 DLL_X1 _10823_ (.D(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__22.cg_i.en_i ),
    .GN(clknet_level_2_1_8164__00543_),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_en ));
 DLL_X1 _10824_ (.D(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__23.cg_i.en_i ),
    .GN(clknet_level_2_1_2146__00543_),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_en ));
 DLL_X1 _10825_ (.D(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__24.cg_i.en_i ),
    .GN(clknet_level_2_1_5155__00543_),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_en ));
 DLL_X1 _10826_ (.D(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__25.cg_i.en_i ),
    .GN(clknet_level_2_1_2146__00543_),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_en ));
 DLL_X1 _10827_ (.D(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__26.cg_i.en_i ),
    .GN(clknet_level_2_1_3149__00543_),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_en ));
 DLL_X1 _10828_ (.D(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__27.cg_i.en_i ),
    .GN(clknet_level_2_1_4152__00543_),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_en ));
 DLL_X1 _10829_ (.D(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__28.cg_i.en_i ),
    .GN(clknet_level_2_1_4152__00543_),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_en ));
 DLL_X1 _10830_ (.D(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__29.cg_i.en_i ),
    .GN(clknet_level_2_1_2146__00543_),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_en ));
 DLL_X1 _10831_ (.D(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__30.cg_i.en_i ),
    .GN(clknet_level_2_1_1143__00543_),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_en ));
 DLL_X1 _10832_ (.D(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__31.cg_i.en_i ),
    .GN(clknet_level_2_1_1143__00543_),
    .Q(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_en ));
 DLH_X1 _10833_ (.D(net320),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[13][0] ));
 DLH_X1 _10834_ (.D(net311),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[13][1] ));
 DLH_X1 _10835_ (.D(net308),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[13][2] ));
 DLH_X1 _10836_ (.D(net302),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[13][3] ));
 DLH_X1 _10837_ (.D(net297),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[13][4] ));
 DLH_X1 _10838_ (.D(net292),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[13][5] ));
 DLH_X1 _10839_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[6] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[13][6] ));
 DLH_X1 _10840_ (.D(net280),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[13][7] ));
 DLH_X1 _10841_ (.D(net321),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[1][0] ));
 DLH_X1 _10842_ (.D(net315),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[1][1] ));
 DLH_X1 _10843_ (.D(net308),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[1][2] ));
 DLH_X1 _10844_ (.D(net302),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[1][3] ));
 DLH_X1 _10845_ (.D(net297),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[1][4] ));
 DLH_X1 _10846_ (.D(net291),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[1][5] ));
 DLH_X1 _10847_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[6] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[1][6] ));
 DLH_X1 _10848_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[7] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[1][7] ));
 DLH_X1 _10849_ (.D(net321),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[26][0] ));
 DLH_X1 _10850_ (.D(net315),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[26][1] ));
 DLH_X1 _10851_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[2] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[26][2] ));
 DLH_X1 _10852_ (.D(net302),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[26][3] ));
 DLH_X1 _10853_ (.D(net297),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[26][4] ));
 DLH_X1 _10854_ (.D(net291),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[26][5] ));
 DLH_X1 _10855_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[6] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[26][6] ));
 DLH_X1 _10856_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[7] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[26][7] ));
 DLH_X1 _10857_ (.D(net321),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[9][0] ));
 DLH_X1 _10858_ (.D(net311),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[9][1] ));
 DLH_X1 _10859_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[2] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[9][2] ));
 DLH_X1 _10860_ (.D(net302),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[9][3] ));
 DLH_X1 _10861_ (.D(net297),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[9][4] ));
 DLH_X1 _10862_ (.D(net292),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[9][5] ));
 DLH_X1 _10863_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[6] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[9][6] ));
 DLH_X1 _10864_ (.D(net280),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[9][7] ));
 DLH_X1 _10865_ (.D(net319),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[0][0] ));
 DLH_X1 _10866_ (.D(net311),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[0][1] ));
 DLH_X1 _10867_ (.D(net306),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[0][2] ));
 DLH_X1 _10868_ (.D(net303),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[0][3] ));
 DLH_X1 _10869_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[4] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[0][4] ));
 DLH_X1 _10870_ (.D(net292),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[0][5] ));
 DLH_X1 _10871_ (.D(net285),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[0][6] ));
 DLH_X1 _10872_ (.D(net280),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[0][7] ));
 DLH_X1 _10873_ (.D(net321),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[20][0] ));
 DLH_X1 _10874_ (.D(net315),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[20][1] ));
 DLH_X1 _10875_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[2] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[20][2] ));
 DLH_X1 _10876_ (.D(net302),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[20][3] ));
 DLH_X1 _10877_ (.D(net297),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[20][4] ));
 DLH_X1 _10878_ (.D(net292),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[20][5] ));
 DLH_X1 _10879_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[6] ),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[20][6] ));
 DLH_X1 _10880_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[7] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[20][7] ));
 DLH_X1 _10881_ (.D(net321),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[2][0] ));
 DLH_X1 _10882_ (.D(net315),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[2][1] ));
 DLH_X1 _10883_ (.D(net308),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[2][2] ));
 DLH_X1 _10884_ (.D(net302),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[2][3] ));
 DLH_X1 _10885_ (.D(net297),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[2][4] ));
 DLH_X1 _10886_ (.D(net291),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[2][5] ));
 DLH_X1 _10887_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[6] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[2][6] ));
 DLH_X1 _10888_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[7] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[2][7] ));
 DLH_X1 _10889_ (.D(net321),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[25][0] ));
 DLH_X1 _10890_ (.D(net311),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[25][1] ));
 DLH_X1 _10891_ (.D(net308),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[25][2] ));
 DLH_X1 _10892_ (.D(net302),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[25][3] ));
 DLH_X1 _10893_ (.D(net297),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[25][4] ));
 DLH_X1 _10894_ (.D(net292),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[25][5] ));
 DLH_X1 _10895_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[6] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[25][6] ));
 DLH_X1 _10896_ (.D(net280),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[25][7] ));
 DLH_X1 _10897_ (.D(net320),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[10][0] ));
 DLH_X1 _10898_ (.D(net310),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[10][1] ));
 DLH_X1 _10899_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[2] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[10][2] ));
 DLH_X1 _10900_ (.D(net302),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[10][3] ));
 DLH_X1 _10901_ (.D(net297),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[10][4] ));
 DLH_X1 _10902_ (.D(net292),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[10][5] ));
 DLH_X1 _10903_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[6] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[10][6] ));
 DLH_X1 _10904_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[7] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[10][7] ));
 DLH_X1 _10905_ (.D(net321),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[3][0] ));
 DLH_X1 _10906_ (.D(net315),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[3][1] ));
 DLH_X1 _10907_ (.D(net308),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[3][2] ));
 DLH_X1 _10908_ (.D(net302),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[3][3] ));
 DLH_X1 _10909_ (.D(net297),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[3][4] ));
 DLH_X1 _10910_ (.D(net291),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[3][5] ));
 DLH_X1 _10911_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[6] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[3][6] ));
 DLH_X1 _10912_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[7] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[3][7] ));
 DLH_X1 _10913_ (.D(net321),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[16][0] ));
 DLH_X1 _10914_ (.D(net315),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[16][1] ));
 DLH_X1 _10915_ (.D(net308),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[16][2] ));
 DLH_X1 _10916_ (.D(net302),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[16][3] ));
 DLH_X1 _10917_ (.D(net297),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[16][4] ));
 DLH_X1 _10918_ (.D(net291),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[16][5] ));
 DLH_X1 _10919_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[6] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[16][6] ));
 DLH_X1 _10920_ (.D(net280),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[16][7] ));
 DLH_X1 _10921_ (.D(net321),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[24][0] ));
 DLH_X1 _10922_ (.D(net315),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[24][1] ));
 DLH_X1 _10923_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[2] ),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[24][2] ));
 DLH_X1 _10924_ (.D(net302),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[24][3] ));
 DLH_X1 _10925_ (.D(net297),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[24][4] ));
 DLH_X1 _10926_ (.D(net291),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[24][5] ));
 DLH_X1 _10927_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[6] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[24][6] ));
 DLH_X1 _10928_ (.D(net280),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[24][7] ));
 DLH_X1 _10929_ (.D(net320),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[4][0] ));
 DLH_X1 _10930_ (.D(net315),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[4][1] ));
 DLH_X1 _10931_ (.D(net308),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[4][2] ));
 DLH_X1 _10932_ (.D(net302),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[4][3] ));
 DLH_X1 _10933_ (.D(net297),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[4][4] ));
 DLH_X1 _10934_ (.D(net292),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[4][5] ));
 DLH_X1 _10935_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[6] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[4][6] ));
 DLH_X1 _10936_ (.D(net280),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[4][7] ));
 DLH_X1 _10937_ (.D(net321),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[15][0] ));
 DLH_X1 _10938_ (.D(net315),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[15][1] ));
 DLH_X1 _10939_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[2] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[15][2] ));
 DLH_X1 _10940_ (.D(net302),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[15][3] ));
 DLH_X1 _10941_ (.D(net297),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[15][4] ));
 DLH_X1 _10942_ (.D(net291),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[15][5] ));
 DLH_X1 _10943_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[6] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[15][6] ));
 DLH_X1 _10944_ (.D(net280),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[15][7] ));
 DLH_X1 _10945_ (.D(net321),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[11][0] ));
 DLH_X1 _10946_ (.D(net315),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[11][1] ));
 DLH_X1 _10947_ (.D(net308),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[11][2] ));
 DLH_X1 _10948_ (.D(net302),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[11][3] ));
 DLH_X1 _10949_ (.D(net297),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[11][4] ));
 DLH_X1 _10950_ (.D(net291),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[11][5] ));
 DLH_X1 _10951_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[6] ),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[11][6] ));
 DLH_X1 _10952_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[7] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[11][7] ));
 DLH_X1 _10953_ (.D(net321),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[5][0] ));
 DLH_X1 _10954_ (.D(net315),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[5][1] ));
 DLH_X1 _10955_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[2] ),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[5][2] ));
 DLH_X1 _10956_ (.D(net302),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[5][3] ));
 DLH_X1 _10957_ (.D(net297),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[5][4] ));
 DLH_X1 _10958_ (.D(net292),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[5][5] ));
 DLH_X1 _10959_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[6] ),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[5][6] ));
 DLH_X1 _10960_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[7] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[5][7] ));
 DLH_X1 _10961_ (.D(net321),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[23][0] ));
 DLH_X1 _10962_ (.D(net315),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[23][1] ));
 DLH_X1 _10963_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[2] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[23][2] ));
 DLH_X1 _10964_ (.D(net302),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[23][3] ));
 DLH_X1 _10965_ (.D(net297),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[23][4] ));
 DLH_X1 _10966_ (.D(net291),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[23][5] ));
 DLH_X1 _10967_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[6] ),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[23][6] ));
 DLH_X1 _10968_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[7] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[23][7] ));
 DLH_X1 _10969_ (.D(net321),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[19][0] ));
 DLH_X1 _10970_ (.D(net315),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[19][1] ));
 DLH_X1 _10971_ (.D(net308),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[19][2] ));
 DLH_X1 _10972_ (.D(net302),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[19][3] ));
 DLH_X1 _10973_ (.D(net297),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[19][4] ));
 DLH_X1 _10974_ (.D(net291),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[19][5] ));
 DLH_X1 _10975_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[6] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[19][6] ));
 DLH_X1 _10976_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[7] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[19][7] ));
 DLH_X1 _10977_ (.D(net321),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[31][0] ));
 DLH_X1 _10978_ (.D(net315),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[31][1] ));
 DLH_X1 _10979_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[2] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[31][2] ));
 DLH_X1 _10980_ (.D(net302),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[31][3] ));
 DLH_X1 _10981_ (.D(net297),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[31][4] ));
 DLH_X1 _10982_ (.D(net291),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[31][5] ));
 DLH_X1 _10983_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[6] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[31][6] ));
 DLH_X1 _10984_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[7] ),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[31][7] ));
 DLH_X1 _10985_ (.D(net320),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[6][0] ));
 DLH_X1 _10986_ (.D(net315),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[6][1] ));
 DLH_X1 _10987_ (.D(net308),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[6][2] ));
 DLH_X1 _10988_ (.D(net302),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[6][3] ));
 DLH_X1 _10989_ (.D(net297),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[6][4] ));
 DLH_X1 _10990_ (.D(net291),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[6][5] ));
 DLH_X1 _10991_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[6] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[6][6] ));
 DLH_X1 _10992_ (.D(net280),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[6][7] ));
 DLH_X1 _10993_ (.D(net321),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[14][0] ));
 DLH_X1 _10994_ (.D(net315),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[14][1] ));
 DLH_X1 _10995_ (.D(net308),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[14][2] ));
 DLH_X1 _10996_ (.D(net302),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[14][3] ));
 DLH_X1 _10997_ (.D(net297),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[14][4] ));
 DLH_X1 _10998_ (.D(net291),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[14][5] ));
 DLH_X1 _10999_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[6] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[14][6] ));
 DLH_X1 _11000_ (.D(net280),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[14][7] ));
 DLH_X1 _11001_ (.D(net321),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[30][0] ));
 DLH_X1 _11002_ (.D(net310),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[30][1] ));
 DLH_X1 _11003_ (.D(net308),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[30][2] ));
 DLH_X1 _11004_ (.D(net302),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[30][3] ));
 DLH_X1 _11005_ (.D(net297),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[30][4] ));
 DLH_X1 _11006_ (.D(net291),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[30][5] ));
 DLH_X1 _11007_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[6] ),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[30][6] ));
 DLH_X1 _11008_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[7] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[30][7] ));
 DLH_X1 _11009_ (.D(net321),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[22][0] ));
 DLH_X1 _11010_ (.D(net315),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[22][1] ));
 DLH_X1 _11011_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[2] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[22][2] ));
 DLH_X1 _11012_ (.D(net302),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[22][3] ));
 DLH_X1 _11013_ (.D(net297),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[22][4] ));
 DLH_X1 _11014_ (.D(net291),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[22][5] ));
 DLH_X1 _11015_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[6] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[22][6] ));
 DLH_X1 _11016_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[7] ),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[22][7] ));
 DLH_X1 _11017_ (.D(net321),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[7][0] ));
 DLH_X1 _11018_ (.D(net315),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[7][1] ));
 DLH_X1 _11019_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[2] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[7][2] ));
 DLH_X1 _11020_ (.D(net302),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[7][3] ));
 DLH_X1 _11021_ (.D(net297),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[7][4] ));
 DLH_X1 _11022_ (.D(net291),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[7][5] ));
 DLH_X1 _11023_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[6] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[7][6] ));
 DLH_X1 _11024_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[7] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[7][7] ));
 DLH_X1 _11025_ (.D(net320),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[29][0] ));
 DLH_X1 _11026_ (.D(net315),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[29][1] ));
 DLH_X1 _11027_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[2] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[29][2] ));
 DLH_X1 _11028_ (.D(net302),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[29][3] ));
 DLH_X1 _11029_ (.D(net297),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[29][4] ));
 DLH_X1 _11030_ (.D(net291),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[29][5] ));
 DLH_X1 _11031_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[6] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[29][6] ));
 DLH_X1 _11032_ (.D(net280),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[29][7] ));
 DLH_X1 _11033_ (.D(net321),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[12][0] ));
 DLH_X1 _11034_ (.D(net315),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[12][1] ));
 DLH_X1 _11035_ (.D(net308),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[12][2] ));
 DLH_X1 _11036_ (.D(net302),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[12][3] ));
 DLH_X1 _11037_ (.D(net297),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[12][4] ));
 DLH_X1 _11038_ (.D(net291),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[12][5] ));
 DLH_X1 _11039_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[6] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[12][6] ));
 DLH_X1 _11040_ (.D(net280),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[12][7] ));
 DLH_X1 _11041_ (.D(net320),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[17][0] ));
 DLH_X1 _11042_ (.D(net315),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[17][1] ));
 DLH_X1 _11043_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[2] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[17][2] ));
 DLH_X1 _11044_ (.D(net302),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[17][3] ));
 DLH_X1 _11045_ (.D(net297),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[17][4] ));
 DLH_X1 _11046_ (.D(net291),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[17][5] ));
 DLH_X1 _11047_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[6] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[17][6] ));
 DLH_X1 _11048_ (.D(net280),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[17][7] ));
 DLH_X1 _11049_ (.D(net321),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[28][0] ));
 DLH_X1 _11050_ (.D(net310),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[28][1] ));
 DLH_X1 _11051_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[2] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[28][2] ));
 DLH_X1 _11052_ (.D(net302),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[28][3] ));
 DLH_X1 _11053_ (.D(net297),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[28][4] ));
 DLH_X1 _11054_ (.D(net291),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[28][5] ));
 DLH_X1 _11055_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[6] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[28][6] ));
 DLH_X1 _11056_ (.D(net280),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[28][7] ));
 DLH_X1 _11057_ (.D(net320),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[8][0] ));
 DLH_X1 _11058_ (.D(net310),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[8][1] ));
 DLH_X1 _11059_ (.D(net308),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[8][2] ));
 DLH_X1 _11060_ (.D(net302),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[8][3] ));
 DLH_X1 _11061_ (.D(net297),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[8][4] ));
 DLH_X1 _11062_ (.D(net291),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[8][5] ));
 DLH_X1 _11063_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[6] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[8][6] ));
 DLH_X1 _11064_ (.D(net280),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[8][7] ));
 DLH_X1 _11065_ (.D(net321),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[21][0] ));
 DLH_X1 _11066_ (.D(net311),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[21][1] ));
 DLH_X1 _11067_ (.D(net308),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[21][2] ));
 DLH_X1 _11068_ (.D(net302),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[21][3] ));
 DLH_X1 _11069_ (.D(net297),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[21][4] ));
 DLH_X1 _11070_ (.D(net291),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[21][5] ));
 DLH_X1 _11071_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[6] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[21][6] ));
 DLH_X1 _11072_ (.D(net280),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[21][7] ));
 DLH_X1 _11073_ (.D(net321),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[27][0] ));
 DLH_X1 _11074_ (.D(net311),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[27][1] ));
 DLH_X1 _11075_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[2] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[27][2] ));
 DLH_X1 _11076_ (.D(net302),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[27][3] ));
 DLH_X1 _11077_ (.D(net297),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[27][4] ));
 DLH_X1 _11078_ (.D(net291),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[27][5] ));
 DLH_X1 _11079_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[6] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[27][6] ));
 DLH_X1 _11080_ (.D(net280),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[27][7] ));
 DLH_X1 _11081_ (.D(net320),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[18][0] ));
 DLH_X1 _11082_ (.D(net315),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[18][1] ));
 DLH_X1 _11083_ (.D(net308),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[18][2] ));
 DLH_X1 _11084_ (.D(net302),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[18][3] ));
 DLH_X1 _11085_ (.D(net297),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[18][4] ));
 DLH_X1 _11086_ (.D(net291),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[18][5] ));
 DLH_X1 _11087_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[6] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[18][6] ));
 DLH_X1 _11088_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[7] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.mem[18][7] ));
 DLL_X1 _11089_ (.D(\lut.gen_sub_units_scm.__11.sub_unit_i.cg_we_global.en_i ),
    .GN(clknet_level_5_1_4320__00532_),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.cg_we_global.clk_en ));
 DLL_X1 _11090_ (.D(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__0.cg_i.en_i ),
    .GN(clknet_level_2_1_5359__00546_),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_en ));
 DLL_X1 _11091_ (.D(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__1.cg_i.en_i ),
    .GN(clknet_level_2_1_2350__00546_),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_en ));
 DLL_X1 _11092_ (.D(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__2.cg_i.en_i ),
    .GN(clknet_level_2_1_3353__00546_),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_en ));
 DLL_X1 _11093_ (.D(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__3.cg_i.en_i ),
    .GN(clknet_level_2_1_7365__00546_),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_en ));
 DLL_X1 _11094_ (.D(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__4.cg_i.en_i ),
    .GN(clknet_level_2_1_5359__00546_),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_en ));
 DLL_X1 _11095_ (.D(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__5.cg_i.en_i ),
    .GN(clknet_level_2_1_8368__00546_),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_en ));
 DLL_X1 _11096_ (.D(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__6.cg_i.en_i ),
    .GN(clknet_level_2_1_1347__00546_),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_en ));
 DLL_X1 _11097_ (.D(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__7.cg_i.en_i ),
    .GN(clknet_level_2_1_8368__00546_),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_en ));
 DLL_X1 _11098_ (.D(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__8.cg_i.en_i ),
    .GN(clknet_level_2_1_2350__00546_),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_en ));
 DLL_X1 _11099_ (.D(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__9.cg_i.en_i ),
    .GN(clknet_level_2_1_6362__00546_),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_en ));
 DLL_X1 _11100_ (.D(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__10.cg_i.en_i ),
    .GN(clknet_level_2_1_8368__00546_),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_en ));
 DLL_X1 _11101_ (.D(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__11.cg_i.en_i ),
    .GN(clknet_level_2_1_3353__00546_),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_en ));
 DLL_X1 _11102_ (.D(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__12.cg_i.en_i ),
    .GN(clknet_level_2_1_3353__00546_),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_en ));
 DLL_X1 _11103_ (.D(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__13.cg_i.en_i ),
    .GN(clknet_level_2_1_5359__00546_),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_en ));
 DLL_X1 _11104_ (.D(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__14.cg_i.en_i ),
    .GN(clknet_level_2_1_3353__00546_),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_en ));
 DLL_X1 _11105_ (.D(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__15.cg_i.en_i ),
    .GN(clknet_level_2_1_1347__00546_),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_en ));
 DLL_X1 _11106_ (.D(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__16.cg_i.en_i ),
    .GN(clknet_level_2_1_1347__00546_),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_en ));
 DLL_X1 _11107_ (.D(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__17.cg_i.en_i ),
    .GN(clknet_level_2_1_6362__00546_),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_en ));
 DLL_X1 _11108_ (.D(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__18.cg_i.en_i ),
    .GN(clknet_level_2_1_4356__00546_),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_en ));
 DLL_X1 _11109_ (.D(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__19.cg_i.en_i ),
    .GN(clknet_level_2_1_2350__00546_),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_en ));
 DLL_X1 _11110_ (.D(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__20.cg_i.en_i ),
    .GN(clknet_level_2_1_8368__00546_),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_en ));
 DLL_X1 _11111_ (.D(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__21.cg_i.en_i ),
    .GN(clknet_level_2_1_6362__00546_),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_en ));
 DLL_X1 _11112_ (.D(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__22.cg_i.en_i ),
    .GN(clknet_level_2_1_3353__00546_),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_en ));
 DLL_X1 _11113_ (.D(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__23.cg_i.en_i ),
    .GN(clknet_level_2_1_4356__00546_),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_en ));
 DLL_X1 _11114_ (.D(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__24.cg_i.en_i ),
    .GN(clknet_level_2_1_2350__00546_),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_en ));
 DLL_X1 _11115_ (.D(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__25.cg_i.en_i ),
    .GN(clknet_level_2_1_6362__00546_),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_en ));
 DLL_X1 _11116_ (.D(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__26.cg_i.en_i ),
    .GN(clknet_level_2_1_5359__00546_),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_en ));
 DLL_X1 _11117_ (.D(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__27.cg_i.en_i ),
    .GN(clknet_level_2_1_5359__00546_),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_en ));
 DLL_X1 _11118_ (.D(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__28.cg_i.en_i ),
    .GN(clknet_level_2_1_1347__00546_),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_en ));
 DLL_X1 _11119_ (.D(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__29.cg_i.en_i ),
    .GN(clknet_level_2_1_1347__00546_),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_en ));
 DLL_X1 _11120_ (.D(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__30.cg_i.en_i ),
    .GN(clknet_level_2_1_3353__00546_),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_en ));
 DLL_X1 _11121_ (.D(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__31.cg_i.en_i ),
    .GN(clknet_level_2_1_4356__00546_),
    .Q(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_en ));
 DLH_X1 _11122_ (.D(net320),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[13][0] ));
 DLH_X1 _11123_ (.D(net311),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[13][1] ));
 DLH_X1 _11124_ (.D(net305),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[13][2] ));
 DLH_X1 _11125_ (.D(net299),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[13][3] ));
 DLH_X1 _11126_ (.D(net294),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[13][4] ));
 DLH_X1 _11127_ (.D(net287),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[13][5] ));
 DLH_X1 _11128_ (.D(net282),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[13][6] ));
 DLH_X1 _11129_ (.D(net275),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[13][7] ));
 DLH_X1 _11130_ (.D(net317),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[1][0] ));
 DLH_X1 _11131_ (.D(net311),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[1][1] ));
 DLH_X1 _11132_ (.D(net305),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[1][2] ));
 DLH_X1 _11133_ (.D(net299),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[1][3] ));
 DLH_X1 _11134_ (.D(net294),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[1][4] ));
 DLH_X1 _11135_ (.D(net287),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[1][5] ));
 DLH_X1 _11136_ (.D(net282),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[1][6] ));
 DLH_X1 _11137_ (.D(net277),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[1][7] ));
 DLH_X1 _11138_ (.D(net317),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[26][0] ));
 DLH_X1 _11139_ (.D(net311),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[26][1] ));
 DLH_X1 _11140_ (.D(net305),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[26][2] ));
 DLH_X1 _11141_ (.D(net299),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[26][3] ));
 DLH_X1 _11142_ (.D(net294),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[26][4] ));
 DLH_X1 _11143_ (.D(net287),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[26][5] ));
 DLH_X1 _11144_ (.D(net282),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[26][6] ));
 DLH_X1 _11145_ (.D(net277),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[26][7] ));
 DLH_X1 _11146_ (.D(net317),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[9][0] ));
 DLH_X1 _11147_ (.D(net311),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[9][1] ));
 DLH_X1 _11148_ (.D(net305),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[9][2] ));
 DLH_X1 _11149_ (.D(net299),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[9][3] ));
 DLH_X1 _11150_ (.D(net294),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[9][4] ));
 DLH_X1 _11151_ (.D(net287),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[9][5] ));
 DLH_X1 _11152_ (.D(net282),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[9][6] ));
 DLH_X1 _11153_ (.D(net277),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[9][7] ));
 DLH_X1 _11154_ (.D(net317),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[0][0] ));
 DLH_X1 _11155_ (.D(net313),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[0][1] ));
 DLH_X1 _11156_ (.D(net305),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[0][2] ));
 DLH_X1 _11157_ (.D(net303),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[0][3] ));
 DLH_X1 _11158_ (.D(net294),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[0][4] ));
 DLH_X1 _11159_ (.D(net287),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[0][5] ));
 DLH_X1 _11160_ (.D(net285),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[0][6] ));
 DLH_X1 _11161_ (.D(net277),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[0][7] ));
 DLH_X1 _11162_ (.D(net320),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[20][0] ));
 DLH_X1 _11163_ (.D(net311),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[20][1] ));
 DLH_X1 _11164_ (.D(net305),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[20][2] ));
 DLH_X1 _11165_ (.D(net299),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[20][3] ));
 DLH_X1 _11166_ (.D(net294),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[20][4] ));
 DLH_X1 _11167_ (.D(net287),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[20][5] ));
 DLH_X1 _11168_ (.D(net282),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[20][6] ));
 DLH_X1 _11169_ (.D(net277),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[20][7] ));
 DLH_X1 _11170_ (.D(net317),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[2][0] ));
 DLH_X1 _11171_ (.D(net311),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[2][1] ));
 DLH_X1 _11172_ (.D(net305),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[2][2] ));
 DLH_X1 _11173_ (.D(net299),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[2][3] ));
 DLH_X1 _11174_ (.D(net294),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[2][4] ));
 DLH_X1 _11175_ (.D(net287),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[2][5] ));
 DLH_X1 _11176_ (.D(net282),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[2][6] ));
 DLH_X1 _11177_ (.D(net277),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[2][7] ));
 DLH_X1 _11178_ (.D(net317),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[25][0] ));
 DLH_X1 _11179_ (.D(net311),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[25][1] ));
 DLH_X1 _11180_ (.D(net305),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[25][2] ));
 DLH_X1 _11181_ (.D(net299),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[25][3] ));
 DLH_X1 _11182_ (.D(net294),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[25][4] ));
 DLH_X1 _11183_ (.D(net287),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[25][5] ));
 DLH_X1 _11184_ (.D(net282),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[25][6] ));
 DLH_X1 _11185_ (.D(net277),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[25][7] ));
 DLH_X1 _11186_ (.D(net320),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[10][0] ));
 DLH_X1 _11187_ (.D(net311),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[10][1] ));
 DLH_X1 _11188_ (.D(net305),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[10][2] ));
 DLH_X1 _11189_ (.D(net299),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[10][3] ));
 DLH_X1 _11190_ (.D(net294),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[10][4] ));
 DLH_X1 _11191_ (.D(net287),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[10][5] ));
 DLH_X1 _11192_ (.D(net282),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[10][6] ));
 DLH_X1 _11193_ (.D(net277),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[10][7] ));
 DLH_X1 _11194_ (.D(net317),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[3][0] ));
 DLH_X1 _11195_ (.D(net311),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[3][1] ));
 DLH_X1 _11196_ (.D(net305),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[3][2] ));
 DLH_X1 _11197_ (.D(net299),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[3][3] ));
 DLH_X1 _11198_ (.D(net294),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[3][4] ));
 DLH_X1 _11199_ (.D(net287),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[3][5] ));
 DLH_X1 _11200_ (.D(net282),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[3][6] ));
 DLH_X1 _11201_ (.D(net277),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[3][7] ));
 DLH_X1 _11202_ (.D(net320),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[16][0] ));
 DLH_X1 _11203_ (.D(net311),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[16][1] ));
 DLH_X1 _11204_ (.D(net305),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[16][2] ));
 DLH_X1 _11205_ (.D(net299),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[16][3] ));
 DLH_X1 _11206_ (.D(net294),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[16][4] ));
 DLH_X1 _11207_ (.D(net287),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[16][5] ));
 DLH_X1 _11208_ (.D(net282),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[16][6] ));
 DLH_X1 _11209_ (.D(net277),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[16][7] ));
 DLH_X1 _11210_ (.D(net320),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[24][0] ));
 DLH_X1 _11211_ (.D(net311),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[24][1] ));
 DLH_X1 _11212_ (.D(net305),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[24][2] ));
 DLH_X1 _11213_ (.D(net299),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[24][3] ));
 DLH_X1 _11214_ (.D(net294),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[24][4] ));
 DLH_X1 _11215_ (.D(net287),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[24][5] ));
 DLH_X1 _11216_ (.D(net282),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[24][6] ));
 DLH_X1 _11217_ (.D(net277),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[24][7] ));
 DLH_X1 _11218_ (.D(net317),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[4][0] ));
 DLH_X1 _11219_ (.D(net311),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[4][1] ));
 DLH_X1 _11220_ (.D(net305),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[4][2] ));
 DLH_X1 _11221_ (.D(net299),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[4][3] ));
 DLH_X1 _11222_ (.D(net294),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[4][4] ));
 DLH_X1 _11223_ (.D(net287),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[4][5] ));
 DLH_X1 _11224_ (.D(net282),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[4][6] ));
 DLH_X1 _11225_ (.D(net277),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[4][7] ));
 DLH_X1 _11226_ (.D(net317),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[15][0] ));
 DLH_X1 _11227_ (.D(net311),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[15][1] ));
 DLH_X1 _11228_ (.D(net305),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[15][2] ));
 DLH_X1 _11229_ (.D(net299),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[15][3] ));
 DLH_X1 _11230_ (.D(net294),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[15][4] ));
 DLH_X1 _11231_ (.D(net287),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[15][5] ));
 DLH_X1 _11232_ (.D(net282),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[15][6] ));
 DLH_X1 _11233_ (.D(net275),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[15][7] ));
 DLH_X1 _11234_ (.D(net317),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[11][0] ));
 DLH_X1 _11235_ (.D(net311),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[11][1] ));
 DLH_X1 _11236_ (.D(net305),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[11][2] ));
 DLH_X1 _11237_ (.D(net299),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[11][3] ));
 DLH_X1 _11238_ (.D(net294),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[11][4] ));
 DLH_X1 _11239_ (.D(net287),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[11][5] ));
 DLH_X1 _11240_ (.D(net282),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[11][6] ));
 DLH_X1 _11241_ (.D(net277),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[11][7] ));
 DLH_X1 _11242_ (.D(net317),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[5][0] ));
 DLH_X1 _11243_ (.D(net311),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[5][1] ));
 DLH_X1 _11244_ (.D(net305),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[5][2] ));
 DLH_X1 _11245_ (.D(net299),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[5][3] ));
 DLH_X1 _11246_ (.D(net294),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[5][4] ));
 DLH_X1 _11247_ (.D(net287),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[5][5] ));
 DLH_X1 _11248_ (.D(net282),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[5][6] ));
 DLH_X1 _11249_ (.D(net277),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[5][7] ));
 DLH_X1 _11250_ (.D(net317),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[23][0] ));
 DLH_X1 _11251_ (.D(net311),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[23][1] ));
 DLH_X1 _11252_ (.D(net305),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[23][2] ));
 DLH_X1 _11253_ (.D(net299),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[23][3] ));
 DLH_X1 _11254_ (.D(net294),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[23][4] ));
 DLH_X1 _11255_ (.D(net287),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[23][5] ));
 DLH_X1 _11256_ (.D(net282),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[23][6] ));
 DLH_X1 _11257_ (.D(net277),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[23][7] ));
 DLH_X1 _11258_ (.D(net317),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[19][0] ));
 DLH_X1 _11259_ (.D(net311),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[19][1] ));
 DLH_X1 _11260_ (.D(net305),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[19][2] ));
 DLH_X1 _11261_ (.D(net299),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[19][3] ));
 DLH_X1 _11262_ (.D(net294),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[19][4] ));
 DLH_X1 _11263_ (.D(net287),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[19][5] ));
 DLH_X1 _11264_ (.D(net282),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[19][6] ));
 DLH_X1 _11265_ (.D(net277),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[19][7] ));
 DLH_X1 _11266_ (.D(net317),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[31][0] ));
 DLH_X1 _11267_ (.D(net311),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[31][1] ));
 DLH_X1 _11268_ (.D(net305),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[31][2] ));
 DLH_X1 _11269_ (.D(net299),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[31][3] ));
 DLH_X1 _11270_ (.D(net294),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[31][4] ));
 DLH_X1 _11271_ (.D(net287),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[31][5] ));
 DLH_X1 _11272_ (.D(net282),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[31][6] ));
 DLH_X1 _11273_ (.D(net277),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[31][7] ));
 DLH_X1 _11274_ (.D(net317),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[6][0] ));
 DLH_X1 _11275_ (.D(net311),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[6][1] ));
 DLH_X1 _11276_ (.D(net305),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[6][2] ));
 DLH_X1 _11277_ (.D(net299),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[6][3] ));
 DLH_X1 _11278_ (.D(net294),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[6][4] ));
 DLH_X1 _11279_ (.D(net287),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[6][5] ));
 DLH_X1 _11280_ (.D(net282),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[6][6] ));
 DLH_X1 _11281_ (.D(net277),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[6][7] ));
 DLH_X1 _11282_ (.D(net320),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[14][0] ));
 DLH_X1 _11283_ (.D(net311),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[14][1] ));
 DLH_X1 _11284_ (.D(net305),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[14][2] ));
 DLH_X1 _11285_ (.D(net299),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[14][3] ));
 DLH_X1 _11286_ (.D(net294),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[14][4] ));
 DLH_X1 _11287_ (.D(net287),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[14][5] ));
 DLH_X1 _11288_ (.D(net282),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[14][6] ));
 DLH_X1 _11289_ (.D(net277),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[14][7] ));
 DLH_X1 _11290_ (.D(net317),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[30][0] ));
 DLH_X1 _11291_ (.D(net311),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[30][1] ));
 DLH_X1 _11292_ (.D(net305),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[30][2] ));
 DLH_X1 _11293_ (.D(net299),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[30][3] ));
 DLH_X1 _11294_ (.D(net294),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[30][4] ));
 DLH_X1 _11295_ (.D(net287),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[30][5] ));
 DLH_X1 _11296_ (.D(net282),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[30][6] ));
 DLH_X1 _11297_ (.D(net277),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[30][7] ));
 DLH_X1 _11298_ (.D(net317),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[22][0] ));
 DLH_X1 _11299_ (.D(net311),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[22][1] ));
 DLH_X1 _11300_ (.D(net305),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[22][2] ));
 DLH_X1 _11301_ (.D(net299),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[22][3] ));
 DLH_X1 _11302_ (.D(net294),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[22][4] ));
 DLH_X1 _11303_ (.D(net287),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[22][5] ));
 DLH_X1 _11304_ (.D(net282),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[22][6] ));
 DLH_X1 _11305_ (.D(net277),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[22][7] ));
 DLH_X1 _11306_ (.D(net317),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[7][0] ));
 DLH_X1 _11307_ (.D(net311),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[7][1] ));
 DLH_X1 _11308_ (.D(net305),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[7][2] ));
 DLH_X1 _11309_ (.D(net299),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[7][3] ));
 DLH_X1 _11310_ (.D(net294),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[7][4] ));
 DLH_X1 _11311_ (.D(net287),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[7][5] ));
 DLH_X1 _11312_ (.D(net282),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[7][6] ));
 DLH_X1 _11313_ (.D(net277),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[7][7] ));
 DLH_X1 _11314_ (.D(net317),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[29][0] ));
 DLH_X1 _11315_ (.D(net311),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[29][1] ));
 DLH_X1 _11316_ (.D(net305),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[29][2] ));
 DLH_X1 _11317_ (.D(net299),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[29][3] ));
 DLH_X1 _11318_ (.D(net294),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[29][4] ));
 DLH_X1 _11319_ (.D(net287),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[29][5] ));
 DLH_X1 _11320_ (.D(net282),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[29][6] ));
 DLH_X1 _11321_ (.D(net277),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[29][7] ));
 DLH_X1 _11322_ (.D(net317),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[12][0] ));
 DLH_X1 _11323_ (.D(net311),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[12][1] ));
 DLH_X1 _11324_ (.D(net305),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[12][2] ));
 DLH_X1 _11325_ (.D(net299),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[12][3] ));
 DLH_X1 _11326_ (.D(net294),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[12][4] ));
 DLH_X1 _11327_ (.D(net287),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[12][5] ));
 DLH_X1 _11328_ (.D(net282),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[12][6] ));
 DLH_X1 _11329_ (.D(net277),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[12][7] ));
 DLH_X1 _11330_ (.D(net317),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[17][0] ));
 DLH_X1 _11331_ (.D(net311),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[17][1] ));
 DLH_X1 _11332_ (.D(net305),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[17][2] ));
 DLH_X1 _11333_ (.D(net299),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[17][3] ));
 DLH_X1 _11334_ (.D(net294),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[17][4] ));
 DLH_X1 _11335_ (.D(net287),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[17][5] ));
 DLH_X1 _11336_ (.D(net282),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[17][6] ));
 DLH_X1 _11337_ (.D(net277),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[17][7] ));
 DLH_X1 _11338_ (.D(net320),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[28][0] ));
 DLH_X1 _11339_ (.D(net311),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[28][1] ));
 DLH_X1 _11340_ (.D(net305),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[28][2] ));
 DLH_X1 _11341_ (.D(net299),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[28][3] ));
 DLH_X1 _11342_ (.D(net294),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[28][4] ));
 DLH_X1 _11343_ (.D(net287),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[28][5] ));
 DLH_X1 _11344_ (.D(net282),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[28][6] ));
 DLH_X1 _11345_ (.D(net277),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[28][7] ));
 DLH_X1 _11346_ (.D(net317),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[8][0] ));
 DLH_X1 _11347_ (.D(net311),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[8][1] ));
 DLH_X1 _11348_ (.D(net305),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[8][2] ));
 DLH_X1 _11349_ (.D(net299),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[8][3] ));
 DLH_X1 _11350_ (.D(net294),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[8][4] ));
 DLH_X1 _11351_ (.D(net287),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[8][5] ));
 DLH_X1 _11352_ (.D(net282),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[8][6] ));
 DLH_X1 _11353_ (.D(net277),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[8][7] ));
 DLH_X1 _11354_ (.D(net317),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[21][0] ));
 DLH_X1 _11355_ (.D(net311),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[21][1] ));
 DLH_X1 _11356_ (.D(net305),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[21][2] ));
 DLH_X1 _11357_ (.D(net299),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[21][3] ));
 DLH_X1 _11358_ (.D(net294),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[21][4] ));
 DLH_X1 _11359_ (.D(net287),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[21][5] ));
 DLH_X1 _11360_ (.D(net282),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[21][6] ));
 DLH_X1 _11361_ (.D(net277),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[21][7] ));
 DLH_X1 _11362_ (.D(net320),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[27][0] ));
 DLH_X1 _11363_ (.D(net311),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[27][1] ));
 DLH_X1 _11364_ (.D(net305),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[27][2] ));
 DLH_X1 _11365_ (.D(net299),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[27][3] ));
 DLH_X1 _11366_ (.D(net294),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[27][4] ));
 DLH_X1 _11367_ (.D(net287),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[27][5] ));
 DLH_X1 _11368_ (.D(net282),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[27][6] ));
 DLH_X1 _11369_ (.D(net277),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[27][7] ));
 DLH_X1 _11370_ (.D(net317),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[18][0] ));
 DLH_X1 _11371_ (.D(net311),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[18][1] ));
 DLH_X1 _11372_ (.D(net305),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[18][2] ));
 DLH_X1 _11373_ (.D(net299),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[18][3] ));
 DLH_X1 _11374_ (.D(net294),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[18][4] ));
 DLH_X1 _11375_ (.D(net287),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[18][5] ));
 DLH_X1 _11376_ (.D(net282),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[18][6] ));
 DLH_X1 _11377_ (.D(net277),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.mem[18][7] ));
 DLL_X1 _11378_ (.D(\lut.gen_sub_units_scm.__10.sub_unit_i.cg_we_global.en_i ),
    .GN(clknet_level_5_1_114__00532_),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.cg_we_global.clk_en ));
 DLL_X1 _11379_ (.D(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__0.cg_i.en_i ),
    .GN(clknet_level_2_1_838__00549_),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_en ));
 DLL_X1 _11380_ (.D(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__1.cg_i.en_i ),
    .GN(clknet_level_2_1_220__00549_),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_en ));
 DLL_X1 _11381_ (.D(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__2.cg_i.en_i ),
    .GN(clknet_level_2_1_117__00549_),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_en ));
 DLL_X1 _11382_ (.D(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__3.cg_i.en_i ),
    .GN(clknet_level_2_1_220__00549_),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_en ));
 DLL_X1 _11383_ (.D(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__4.cg_i.en_i ),
    .GN(clknet_level_2_1_117__00549_),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_en ));
 DLL_X1 _11384_ (.D(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__5.cg_i.en_i ),
    .GN(clknet_level_2_1_323__00549_),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_en ));
 DLL_X1 _11385_ (.D(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__6.cg_i.en_i ),
    .GN(clknet_level_2_1_426__00549_),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_en ));
 DLL_X1 _11386_ (.D(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__7.cg_i.en_i ),
    .GN(clknet_level_2_1_117__00549_),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_en ));
 DLL_X1 _11387_ (.D(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__8.cg_i.en_i ),
    .GN(clknet_level_2_1_735__00549_),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_en ));
 DLL_X1 _11388_ (.D(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__9.cg_i.en_i ),
    .GN(clknet_level_2_1_529__00549_),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_en ));
 DLL_X1 _11389_ (.D(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__10.cg_i.en_i ),
    .GN(clknet_level_2_1_323__00549_),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_en ));
 DLL_X1 _11390_ (.D(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__11.cg_i.en_i ),
    .GN(clknet_level_2_1_323__00549_),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_en ));
 DLL_X1 _11391_ (.D(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__12.cg_i.en_i ),
    .GN(clknet_level_2_1_220__00549_),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_en ));
 DLL_X1 _11392_ (.D(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__13.cg_i.en_i ),
    .GN(clknet_level_2_1_632__00549_),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_en ));
 DLL_X1 _11393_ (.D(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__14.cg_i.en_i ),
    .GN(clknet_level_2_1_529__00549_),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_en ));
 DLL_X1 _11394_ (.D(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__15.cg_i.en_i ),
    .GN(clknet_level_2_1_220__00549_),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_en ));
 DLL_X1 _11395_ (.D(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__16.cg_i.en_i ),
    .GN(clknet_level_2_1_632__00549_),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_en ));
 DLL_X1 _11396_ (.D(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__17.cg_i.en_i ),
    .GN(clknet_level_2_1_323__00549_),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_en ));
 DLL_X1 _11397_ (.D(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__18.cg_i.en_i ),
    .GN(clknet_level_2_1_632__00549_),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_en ));
 DLL_X1 _11398_ (.D(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__19.cg_i.en_i ),
    .GN(clknet_level_2_1_220__00549_),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_en ));
 DLL_X1 _11399_ (.D(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__20.cg_i.en_i ),
    .GN(clknet_level_2_1_632__00549_),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_en ));
 DLL_X1 _11400_ (.D(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__21.cg_i.en_i ),
    .GN(clknet_level_2_1_426__00549_),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_en ));
 DLL_X1 _11401_ (.D(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__22.cg_i.en_i ),
    .GN(clknet_level_2_1_838__00549_),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_en ));
 DLL_X1 _11402_ (.D(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__23.cg_i.en_i ),
    .GN(clknet_level_2_1_426__00549_),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_en ));
 DLL_X1 _11403_ (.D(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__24.cg_i.en_i ),
    .GN(clknet_level_2_1_529__00549_),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_en ));
 DLL_X1 _11404_ (.D(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__25.cg_i.en_i ),
    .GN(clknet_level_2_1_735__00549_),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_en ));
 DLL_X1 _11405_ (.D(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__26.cg_i.en_i ),
    .GN(clknet_level_2_1_117__00549_),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_en ));
 DLL_X1 _11406_ (.D(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__27.cg_i.en_i ),
    .GN(clknet_level_2_1_735__00549_),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_en ));
 DLL_X1 _11407_ (.D(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__28.cg_i.en_i ),
    .GN(clknet_level_2_1_838__00549_),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_en ));
 DLL_X1 _11408_ (.D(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__29.cg_i.en_i ),
    .GN(clknet_level_2_1_117__00549_),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_en ));
 DLL_X1 _11409_ (.D(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__30.cg_i.en_i ),
    .GN(clknet_level_2_1_426__00549_),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_en ));
 DLL_X1 _11410_ (.D(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__31.cg_i.en_i ),
    .GN(clknet_level_2_1_117__00549_),
    .Q(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_en ));
 DLH_X1 _11411_ (.D(net319),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[13][0] ));
 DLH_X1 _11412_ (.D(net312),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[13][1] ));
 DLH_X1 _11413_ (.D(net304),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[13][2] ));
 DLH_X1 _11414_ (.D(net298),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[13][3] ));
 DLH_X1 _11415_ (.D(net295),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[13][4] ));
 DLH_X1 _11416_ (.D(net289),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[13][5] ));
 DLH_X1 _11417_ (.D(net281),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[13][6] ));
 DLH_X1 _11418_ (.D(net279),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[13][7] ));
 DLH_X1 _11419_ (.D(net319),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[1][0] ));
 DLH_X1 _11420_ (.D(net312),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[1][1] ));
 DLH_X1 _11421_ (.D(net304),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[1][2] ));
 DLH_X1 _11422_ (.D(net298),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[1][3] ));
 DLH_X1 _11423_ (.D(net295),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[1][4] ));
 DLH_X1 _11424_ (.D(net289),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[1][5] ));
 DLH_X1 _11425_ (.D(net281),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[1][6] ));
 DLH_X1 _11426_ (.D(net279),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[1][7] ));
 DLH_X1 _11427_ (.D(net319),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[26][0] ));
 DLH_X1 _11428_ (.D(net312),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[26][1] ));
 DLH_X1 _11429_ (.D(net304),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[26][2] ));
 DLH_X1 _11430_ (.D(net298),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[26][3] ));
 DLH_X1 _11431_ (.D(net295),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[26][4] ));
 DLH_X1 _11432_ (.D(net289),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[26][5] ));
 DLH_X1 _11433_ (.D(net281),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[26][6] ));
 DLH_X1 _11434_ (.D(net279),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[26][7] ));
 DLH_X1 _11435_ (.D(net319),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[9][0] ));
 DLH_X1 _11436_ (.D(net312),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[9][1] ));
 DLH_X1 _11437_ (.D(net304),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[9][2] ));
 DLH_X1 _11438_ (.D(net298),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[9][3] ));
 DLH_X1 _11439_ (.D(net295),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[9][4] ));
 DLH_X1 _11440_ (.D(net289),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[9][5] ));
 DLH_X1 _11441_ (.D(net281),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[9][6] ));
 DLH_X1 _11442_ (.D(net279),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[9][7] ));
 DLH_X1 _11443_ (.D(net319),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[0][0] ));
 DLH_X1 _11444_ (.D(net312),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[0][1] ));
 DLH_X1 _11445_ (.D(net304),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[0][2] ));
 DLH_X1 _11446_ (.D(net298),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[0][3] ));
 DLH_X1 _11447_ (.D(net295),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[0][4] ));
 DLH_X1 _11448_ (.D(net292),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[0][5] ));
 DLH_X1 _11449_ (.D(net285),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[0][6] ));
 DLH_X1 _11450_ (.D(net277),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[0][7] ));
 DLH_X1 _11451_ (.D(net319),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[20][0] ));
 DLH_X1 _11452_ (.D(net312),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[20][1] ));
 DLH_X1 _11453_ (.D(net304),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[20][2] ));
 DLH_X1 _11454_ (.D(net298),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[20][3] ));
 DLH_X1 _11455_ (.D(net296),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[20][4] ));
 DLH_X1 _11456_ (.D(net289),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[20][5] ));
 DLH_X1 _11457_ (.D(net281),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[20][6] ));
 DLH_X1 _11458_ (.D(net279),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[20][7] ));
 DLH_X1 _11459_ (.D(net319),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[2][0] ));
 DLH_X1 _11460_ (.D(net312),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[2][1] ));
 DLH_X1 _11461_ (.D(net304),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[2][2] ));
 DLH_X1 _11462_ (.D(net298),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[2][3] ));
 DLH_X1 _11463_ (.D(net296),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[2][4] ));
 DLH_X1 _11464_ (.D(net289),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[2][5] ));
 DLH_X1 _11465_ (.D(net281),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[2][6] ));
 DLH_X1 _11466_ (.D(net279),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[2][7] ));
 DLH_X1 _11467_ (.D(net319),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[25][0] ));
 DLH_X1 _11468_ (.D(net312),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[25][1] ));
 DLH_X1 _11469_ (.D(net304),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[25][2] ));
 DLH_X1 _11470_ (.D(net298),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[25][3] ));
 DLH_X1 _11471_ (.D(net295),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[25][4] ));
 DLH_X1 _11472_ (.D(net289),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[25][5] ));
 DLH_X1 _11473_ (.D(net281),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[25][6] ));
 DLH_X1 _11474_ (.D(net279),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[25][7] ));
 DLH_X1 _11475_ (.D(net319),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[10][0] ));
 DLH_X1 _11476_ (.D(net312),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[10][1] ));
 DLH_X1 _11477_ (.D(net304),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[10][2] ));
 DLH_X1 _11478_ (.D(net298),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[10][3] ));
 DLH_X1 _11479_ (.D(net295),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[10][4] ));
 DLH_X1 _11480_ (.D(net289),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[10][5] ));
 DLH_X1 _11481_ (.D(net281),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[10][6] ));
 DLH_X1 _11482_ (.D(net279),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[10][7] ));
 DLH_X1 _11483_ (.D(net316),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[3][0] ));
 DLH_X1 _11484_ (.D(net312),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[3][1] ));
 DLH_X1 _11485_ (.D(net304),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[3][2] ));
 DLH_X1 _11486_ (.D(net298),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[3][3] ));
 DLH_X1 _11487_ (.D(net295),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[3][4] ));
 DLH_X1 _11488_ (.D(net289),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[3][5] ));
 DLH_X1 _11489_ (.D(net281),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[3][6] ));
 DLH_X1 _11490_ (.D(net279),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[3][7] ));
 DLH_X1 _11491_ (.D(net319),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[16][0] ));
 DLH_X1 _11492_ (.D(net312),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[16][1] ));
 DLH_X1 _11493_ (.D(net304),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[16][2] ));
 DLH_X1 _11494_ (.D(net298),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[16][3] ));
 DLH_X1 _11495_ (.D(net295),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[16][4] ));
 DLH_X1 _11496_ (.D(net289),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[16][5] ));
 DLH_X1 _11497_ (.D(net281),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[16][6] ));
 DLH_X1 _11498_ (.D(net279),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[16][7] ));
 DLH_X1 _11499_ (.D(net319),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[24][0] ));
 DLH_X1 _11500_ (.D(net312),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[24][1] ));
 DLH_X1 _11501_ (.D(net304),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[24][2] ));
 DLH_X1 _11502_ (.D(net298),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[24][3] ));
 DLH_X1 _11503_ (.D(net295),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[24][4] ));
 DLH_X1 _11504_ (.D(net289),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[24][5] ));
 DLH_X1 _11505_ (.D(net281),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[24][6] ));
 DLH_X1 _11506_ (.D(net279),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[24][7] ));
 DLH_X1 _11507_ (.D(net316),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[4][0] ));
 DLH_X1 _11508_ (.D(net312),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[4][1] ));
 DLH_X1 _11509_ (.D(net304),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[4][2] ));
 DLH_X1 _11510_ (.D(net298),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[4][3] ));
 DLH_X1 _11511_ (.D(net295),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[4][4] ));
 DLH_X1 _11512_ (.D(net289),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[4][5] ));
 DLH_X1 _11513_ (.D(net281),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[4][6] ));
 DLH_X1 _11514_ (.D(net279),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[4][7] ));
 DLH_X1 _11515_ (.D(net319),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[15][0] ));
 DLH_X1 _11516_ (.D(net312),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[15][1] ));
 DLH_X1 _11517_ (.D(net304),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[15][2] ));
 DLH_X1 _11518_ (.D(net298),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[15][3] ));
 DLH_X1 _11519_ (.D(net295),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[15][4] ));
 DLH_X1 _11520_ (.D(net289),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[15][5] ));
 DLH_X1 _11521_ (.D(net281),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[15][6] ));
 DLH_X1 _11522_ (.D(net279),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[15][7] ));
 DLH_X1 _11523_ (.D(net319),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[11][0] ));
 DLH_X1 _11524_ (.D(net312),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[11][1] ));
 DLH_X1 _11525_ (.D(net304),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[11][2] ));
 DLH_X1 _11526_ (.D(net298),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[11][3] ));
 DLH_X1 _11527_ (.D(net295),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[11][4] ));
 DLH_X1 _11528_ (.D(net289),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[11][5] ));
 DLH_X1 _11529_ (.D(net281),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[11][6] ));
 DLH_X1 _11530_ (.D(net279),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[11][7] ));
 DLH_X1 _11531_ (.D(net319),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[5][0] ));
 DLH_X1 _11532_ (.D(net312),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[5][1] ));
 DLH_X1 _11533_ (.D(net304),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[5][2] ));
 DLH_X1 _11534_ (.D(net298),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[5][3] ));
 DLH_X1 _11535_ (.D(net296),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[5][4] ));
 DLH_X1 _11536_ (.D(net289),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[5][5] ));
 DLH_X1 _11537_ (.D(net281),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[5][6] ));
 DLH_X1 _11538_ (.D(net279),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[5][7] ));
 DLH_X1 _11539_ (.D(net316),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[23][0] ));
 DLH_X1 _11540_ (.D(net312),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[23][1] ));
 DLH_X1 _11541_ (.D(net304),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[23][2] ));
 DLH_X1 _11542_ (.D(net298),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[23][3] ));
 DLH_X1 _11543_ (.D(net296),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[23][4] ));
 DLH_X1 _11544_ (.D(net289),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[23][5] ));
 DLH_X1 _11545_ (.D(net281),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[23][6] ));
 DLH_X1 _11546_ (.D(net279),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[23][7] ));
 DLH_X1 _11547_ (.D(net319),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[19][0] ));
 DLH_X1 _11548_ (.D(net312),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[19][1] ));
 DLH_X1 _11549_ (.D(net304),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[19][2] ));
 DLH_X1 _11550_ (.D(net298),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[19][3] ));
 DLH_X1 _11551_ (.D(net296),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[19][4] ));
 DLH_X1 _11552_ (.D(net289),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[19][5] ));
 DLH_X1 _11553_ (.D(net281),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[19][6] ));
 DLH_X1 _11554_ (.D(net279),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[19][7] ));
 DLH_X1 _11555_ (.D(net316),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[31][0] ));
 DLH_X1 _11556_ (.D(net312),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[31][1] ));
 DLH_X1 _11557_ (.D(net304),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[31][2] ));
 DLH_X1 _11558_ (.D(net298),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[31][3] ));
 DLH_X1 _11559_ (.D(net295),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[31][4] ));
 DLH_X1 _11560_ (.D(net289),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[31][5] ));
 DLH_X1 _11561_ (.D(net281),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[31][6] ));
 DLH_X1 _11562_ (.D(net279),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[31][7] ));
 DLH_X1 _11563_ (.D(net319),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[6][0] ));
 DLH_X1 _11564_ (.D(net312),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[6][1] ));
 DLH_X1 _11565_ (.D(net304),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[6][2] ));
 DLH_X1 _11566_ (.D(net298),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[6][3] ));
 DLH_X1 _11567_ (.D(net296),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[6][4] ));
 DLH_X1 _11568_ (.D(net289),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[6][5] ));
 DLH_X1 _11569_ (.D(net281),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[6][6] ));
 DLH_X1 _11570_ (.D(net279),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[6][7] ));
 DLH_X1 _11571_ (.D(net319),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[14][0] ));
 DLH_X1 _11572_ (.D(net312),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[14][1] ));
 DLH_X1 _11573_ (.D(net304),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[14][2] ));
 DLH_X1 _11574_ (.D(net298),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[14][3] ));
 DLH_X1 _11575_ (.D(net295),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[14][4] ));
 DLH_X1 _11576_ (.D(net289),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[14][5] ));
 DLH_X1 _11577_ (.D(net281),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[14][6] ));
 DLH_X1 _11578_ (.D(net279),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[14][7] ));
 DLH_X1 _11579_ (.D(net319),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[30][0] ));
 DLH_X1 _11580_ (.D(net312),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[30][1] ));
 DLH_X1 _11581_ (.D(net304),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[30][2] ));
 DLH_X1 _11582_ (.D(net298),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[30][3] ));
 DLH_X1 _11583_ (.D(net296),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[30][4] ));
 DLH_X1 _11584_ (.D(net289),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[30][5] ));
 DLH_X1 _11585_ (.D(net281),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[30][6] ));
 DLH_X1 _11586_ (.D(net279),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[30][7] ));
 DLH_X1 _11587_ (.D(net319),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[22][0] ));
 DLH_X1 _11588_ (.D(net312),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[22][1] ));
 DLH_X1 _11589_ (.D(net304),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[22][2] ));
 DLH_X1 _11590_ (.D(net298),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[22][3] ));
 DLH_X1 _11591_ (.D(net296),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[22][4] ));
 DLH_X1 _11592_ (.D(net289),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[22][5] ));
 DLH_X1 _11593_ (.D(net281),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[22][6] ));
 DLH_X1 _11594_ (.D(net279),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[22][7] ));
 DLH_X1 _11595_ (.D(net316),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[7][0] ));
 DLH_X1 _11596_ (.D(net312),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[7][1] ));
 DLH_X1 _11597_ (.D(net304),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[7][2] ));
 DLH_X1 _11598_ (.D(net298),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[7][3] ));
 DLH_X1 _11599_ (.D(net295),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[7][4] ));
 DLH_X1 _11600_ (.D(net289),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[7][5] ));
 DLH_X1 _11601_ (.D(net281),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[7][6] ));
 DLH_X1 _11602_ (.D(net279),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[7][7] ));
 DLH_X1 _11603_ (.D(net319),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[29][0] ));
 DLH_X1 _11604_ (.D(net312),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[29][1] ));
 DLH_X1 _11605_ (.D(net304),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[29][2] ));
 DLH_X1 _11606_ (.D(net298),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[29][3] ));
 DLH_X1 _11607_ (.D(net295),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[29][4] ));
 DLH_X1 _11608_ (.D(net289),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[29][5] ));
 DLH_X1 _11609_ (.D(net281),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[29][6] ));
 DLH_X1 _11610_ (.D(net279),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[29][7] ));
 DLH_X1 _11611_ (.D(net319),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[12][0] ));
 DLH_X1 _11612_ (.D(net312),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[12][1] ));
 DLH_X1 _11613_ (.D(net304),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[12][2] ));
 DLH_X1 _11614_ (.D(net298),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[12][3] ));
 DLH_X1 _11615_ (.D(net295),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[12][4] ));
 DLH_X1 _11616_ (.D(net289),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[12][5] ));
 DLH_X1 _11617_ (.D(net281),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[12][6] ));
 DLH_X1 _11618_ (.D(net279),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[12][7] ));
 DLH_X1 _11619_ (.D(net319),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[17][0] ));
 DLH_X1 _11620_ (.D(net312),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[17][1] ));
 DLH_X1 _11621_ (.D(net304),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[17][2] ));
 DLH_X1 _11622_ (.D(net298),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[17][3] ));
 DLH_X1 _11623_ (.D(net295),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[17][4] ));
 DLH_X1 _11624_ (.D(net289),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[17][5] ));
 DLH_X1 _11625_ (.D(net281),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[17][6] ));
 DLH_X1 _11626_ (.D(net279),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[17][7] ));
 DLH_X1 _11627_ (.D(net319),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[28][0] ));
 DLH_X1 _11628_ (.D(net312),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[28][1] ));
 DLH_X1 _11629_ (.D(net304),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[28][2] ));
 DLH_X1 _11630_ (.D(net298),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[28][3] ));
 DLH_X1 _11631_ (.D(net295),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[28][4] ));
 DLH_X1 _11632_ (.D(net289),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[28][5] ));
 DLH_X1 _11633_ (.D(net281),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[28][6] ));
 DLH_X1 _11634_ (.D(net279),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[28][7] ));
 DLH_X1 _11635_ (.D(net319),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[8][0] ));
 DLH_X1 _11636_ (.D(net312),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[8][1] ));
 DLH_X1 _11637_ (.D(net304),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[8][2] ));
 DLH_X1 _11638_ (.D(net298),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[8][3] ));
 DLH_X1 _11639_ (.D(net295),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[8][4] ));
 DLH_X1 _11640_ (.D(net289),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[8][5] ));
 DLH_X1 _11641_ (.D(net281),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[8][6] ));
 DLH_X1 _11642_ (.D(net279),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[8][7] ));
 DLH_X1 _11643_ (.D(net319),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[21][0] ));
 DLH_X1 _11644_ (.D(net312),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[21][1] ));
 DLH_X1 _11645_ (.D(net304),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[21][2] ));
 DLH_X1 _11646_ (.D(net298),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[21][3] ));
 DLH_X1 _11647_ (.D(net295),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[21][4] ));
 DLH_X1 _11648_ (.D(net289),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[21][5] ));
 DLH_X1 _11649_ (.D(net281),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[21][6] ));
 DLH_X1 _11650_ (.D(net279),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[21][7] ));
 DLH_X1 _11651_ (.D(net319),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[27][0] ));
 DLH_X1 _11652_ (.D(net312),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[27][1] ));
 DLH_X1 _11653_ (.D(net304),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[27][2] ));
 DLH_X1 _11654_ (.D(net298),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[27][3] ));
 DLH_X1 _11655_ (.D(net295),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[27][4] ));
 DLH_X1 _11656_ (.D(net289),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[27][5] ));
 DLH_X1 _11657_ (.D(net281),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[27][6] ));
 DLH_X1 _11658_ (.D(net279),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[27][7] ));
 DLH_X1 _11659_ (.D(net319),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[18][0] ));
 DLH_X1 _11660_ (.D(net312),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[18][1] ));
 DLH_X1 _11661_ (.D(net304),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[18][2] ));
 DLH_X1 _11662_ (.D(net298),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[18][3] ));
 DLH_X1 _11663_ (.D(net295),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[18][4] ));
 DLH_X1 _11664_ (.D(net289),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[18][5] ));
 DLH_X1 _11665_ (.D(net281),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[18][6] ));
 DLH_X1 _11666_ (.D(net279),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.mem[18][7] ));
 DLL_X1 _11667_ (.D(\lut.gen_sub_units_scm.__9.sub_unit_i.cg_we_global.en_i ),
    .GN(clknet_level_5_1_2116__00532_),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.cg_we_global.clk_en ));
 DLL_X1 _11668_ (.D(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__0.cg_i.en_i ),
    .GN(clknet_level_2_1_7185__00552_),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_en ));
 DLL_X1 _11669_ (.D(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__1.cg_i.en_i ),
    .GN(clknet_level_2_1_3173__00552_),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_en ));
 DLL_X1 _11670_ (.D(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__2.cg_i.en_i ),
    .GN(clknet_level_2_1_8188__00552_),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_en ));
 DLL_X1 _11671_ (.D(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__3.cg_i.en_i ),
    .GN(clknet_level_2_1_3173__00552_),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_en ));
 DLL_X1 _11672_ (.D(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__4.cg_i.en_i ),
    .GN(clknet_level_2_1_2170__00552_),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_en ));
 DLL_X1 _11673_ (.D(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__5.cg_i.en_i ),
    .GN(clknet_level_2_1_4176__00552_),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_en ));
 DLL_X1 _11674_ (.D(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__6.cg_i.en_i ),
    .GN(clknet_level_2_1_6182__00552_),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_en ));
 DLL_X1 _11675_ (.D(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__7.cg_i.en_i ),
    .GN(clknet_level_2_1_3173__00552_),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_en ));
 DLL_X1 _11676_ (.D(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__8.cg_i.en_i ),
    .GN(clknet_level_2_1_1167__00552_),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_en ));
 DLL_X1 _11677_ (.D(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__9.cg_i.en_i ),
    .GN(clknet_level_2_1_6182__00552_),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_en ));
 DLL_X1 _11678_ (.D(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__10.cg_i.en_i ),
    .GN(clknet_level_2_1_2170__00552_),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_en ));
 DLL_X1 _11679_ (.D(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__11.cg_i.en_i ),
    .GN(clknet_level_2_1_8188__00552_),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_en ));
 DLL_X1 _11680_ (.D(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__12.cg_i.en_i ),
    .GN(clknet_level_2_1_8188__00552_),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_en ));
 DLL_X1 _11681_ (.D(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__13.cg_i.en_i ),
    .GN(clknet_level_2_1_5179__00552_),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_en ));
 DLL_X1 _11682_ (.D(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__14.cg_i.en_i ),
    .GN(clknet_level_2_1_7185__00552_),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_en ));
 DLL_X1 _11683_ (.D(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__15.cg_i.en_i ),
    .GN(clknet_level_2_1_3173__00552_),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_en ));
 DLL_X1 _11684_ (.D(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__16.cg_i.en_i ),
    .GN(clknet_level_2_1_2170__00552_),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_en ));
 DLL_X1 _11685_ (.D(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__17.cg_i.en_i ),
    .GN(clknet_level_2_1_7185__00552_),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_en ));
 DLL_X1 _11686_ (.D(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__18.cg_i.en_i ),
    .GN(clknet_level_2_1_8188__00552_),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_en ));
 DLL_X1 _11687_ (.D(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__19.cg_i.en_i ),
    .GN(clknet_level_2_1_5179__00552_),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_en ));
 DLL_X1 _11688_ (.D(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__20.cg_i.en_i ),
    .GN(clknet_level_2_1_5179__00552_),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_en ));
 DLL_X1 _11689_ (.D(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__21.cg_i.en_i ),
    .GN(clknet_level_2_1_8188__00552_),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_en ));
 DLL_X1 _11690_ (.D(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__22.cg_i.en_i ),
    .GN(clknet_level_2_1_6182__00552_),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_en ));
 DLL_X1 _11691_ (.D(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__23.cg_i.en_i ),
    .GN(clknet_level_2_1_2170__00552_),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_en ));
 DLL_X1 _11692_ (.D(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__24.cg_i.en_i ),
    .GN(clknet_level_2_1_3173__00552_),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_en ));
 DLL_X1 _11693_ (.D(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__25.cg_i.en_i ),
    .GN(clknet_level_2_1_6182__00552_),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_en ));
 DLL_X1 _11694_ (.D(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__26.cg_i.en_i ),
    .GN(clknet_level_2_1_6182__00552_),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_en ));
 DLL_X1 _11695_ (.D(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__27.cg_i.en_i ),
    .GN(clknet_level_2_1_4176__00552_),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_en ));
 DLL_X1 _11696_ (.D(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__28.cg_i.en_i ),
    .GN(clknet_level_2_1_4176__00552_),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_en ));
 DLL_X1 _11697_ (.D(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__29.cg_i.en_i ),
    .GN(clknet_level_2_1_4176__00552_),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_en ));
 DLL_X1 _11698_ (.D(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__30.cg_i.en_i ),
    .GN(clknet_level_2_1_5179__00552_),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_en ));
 DLL_X1 _11699_ (.D(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__31.cg_i.en_i ),
    .GN(clknet_level_2_1_1167__00552_),
    .Q(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_en ));
 DLH_X1 _11700_ (.D(net316),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[13][0] ));
 DLH_X1 _11701_ (.D(net313),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[13][1] ));
 DLH_X1 _11702_ (.D(net304),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[13][2] ));
 DLH_X1 _11703_ (.D(net298),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[13][3] ));
 DLH_X1 _11704_ (.D(net294),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[13][4] ));
 DLH_X1 _11705_ (.D(net288),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[13][5] ));
 DLH_X1 _11706_ (.D(net282),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[13][6] ));
 DLH_X1 _11707_ (.D(net276),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[13][7] ));
 DLH_X1 _11708_ (.D(net316),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[1][0] ));
 DLH_X1 _11709_ (.D(net313),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[1][1] ));
 DLH_X1 _11710_ (.D(net304),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[1][2] ));
 DLH_X1 _11711_ (.D(net298),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[1][3] ));
 DLH_X1 _11712_ (.D(net294),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[1][4] ));
 DLH_X1 _11713_ (.D(net288),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[1][5] ));
 DLH_X1 _11714_ (.D(net282),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[1][6] ));
 DLH_X1 _11715_ (.D(net276),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[1][7] ));
 DLH_X1 _11716_ (.D(net316),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[26][0] ));
 DLH_X1 _11717_ (.D(net313),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[26][1] ));
 DLH_X1 _11718_ (.D(net305),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[26][2] ));
 DLH_X1 _11719_ (.D(net299),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[26][3] ));
 DLH_X1 _11720_ (.D(net294),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[26][4] ));
 DLH_X1 _11721_ (.D(net288),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[26][5] ));
 DLH_X1 _11722_ (.D(net282),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[26][6] ));
 DLH_X1 _11723_ (.D(net276),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[26][7] ));
 DLH_X1 _11724_ (.D(net316),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[9][0] ));
 DLH_X1 _11725_ (.D(net312),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[9][1] ));
 DLH_X1 _11726_ (.D(net305),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[9][2] ));
 DLH_X1 _11727_ (.D(net299),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[9][3] ));
 DLH_X1 _11728_ (.D(net294),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[9][4] ));
 DLH_X1 _11729_ (.D(net288),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[9][5] ));
 DLH_X1 _11730_ (.D(net282),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[9][6] ));
 DLH_X1 _11731_ (.D(net276),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[9][7] ));
 DLH_X1 _11732_ (.D(net316),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[0][0] ));
 DLH_X1 _11733_ (.D(net313),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[0][1] ));
 DLH_X1 _11734_ (.D(net306),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[0][2] ));
 DLH_X1 _11735_ (.D(net298),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[0][3] ));
 DLH_X1 _11736_ (.D(net295),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[0][4] ));
 DLH_X1 _11737_ (.D(net288),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[0][5] ));
 DLH_X1 _11738_ (.D(net282),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[0][6] ));
 DLH_X1 _11739_ (.D(net279),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[0][7] ));
 DLH_X1 _11740_ (.D(net316),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[20][0] ));
 DLH_X1 _11741_ (.D(net313),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[20][1] ));
 DLH_X1 _11742_ (.D(net304),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[20][2] ));
 DLH_X1 _11743_ (.D(net299),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[20][3] ));
 DLH_X1 _11744_ (.D(net294),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[20][4] ));
 DLH_X1 _11745_ (.D(net288),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[20][5] ));
 DLH_X1 _11746_ (.D(net282),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[20][6] ));
 DLH_X1 _11747_ (.D(net276),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[20][7] ));
 DLH_X1 _11748_ (.D(net316),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[2][0] ));
 DLH_X1 _11749_ (.D(net313),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[2][1] ));
 DLH_X1 _11750_ (.D(net305),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[2][2] ));
 DLH_X1 _11751_ (.D(net298),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[2][3] ));
 DLH_X1 _11752_ (.D(net294),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[2][4] ));
 DLH_X1 _11753_ (.D(net288),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[2][5] ));
 DLH_X1 _11754_ (.D(net282),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[2][6] ));
 DLH_X1 _11755_ (.D(net276),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[2][7] ));
 DLH_X1 _11756_ (.D(net316),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[25][0] ));
 DLH_X1 _11757_ (.D(net313),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[25][1] ));
 DLH_X1 _11758_ (.D(net304),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[25][2] ));
 DLH_X1 _11759_ (.D(net298),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[25][3] ));
 DLH_X1 _11760_ (.D(net294),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[25][4] ));
 DLH_X1 _11761_ (.D(net288),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[25][5] ));
 DLH_X1 _11762_ (.D(net282),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[25][6] ));
 DLH_X1 _11763_ (.D(net276),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[25][7] ));
 DLH_X1 _11764_ (.D(net316),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[10][0] ));
 DLH_X1 _11765_ (.D(net312),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[10][1] ));
 DLH_X1 _11766_ (.D(net304),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[10][2] ));
 DLH_X1 _11767_ (.D(net299),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[10][3] ));
 DLH_X1 _11768_ (.D(net294),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[10][4] ));
 DLH_X1 _11769_ (.D(net288),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[10][5] ));
 DLH_X1 _11770_ (.D(net282),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[10][6] ));
 DLH_X1 _11771_ (.D(net276),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[10][7] ));
 DLH_X1 _11772_ (.D(net316),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[3][0] ));
 DLH_X1 _11773_ (.D(net313),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[3][1] ));
 DLH_X1 _11774_ (.D(net305),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[3][2] ));
 DLH_X1 _11775_ (.D(net299),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[3][3] ));
 DLH_X1 _11776_ (.D(net294),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[3][4] ));
 DLH_X1 _11777_ (.D(net288),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[3][5] ));
 DLH_X1 _11778_ (.D(net282),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[3][6] ));
 DLH_X1 _11779_ (.D(net276),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[3][7] ));
 DLH_X1 _11780_ (.D(net316),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[16][0] ));
 DLH_X1 _11781_ (.D(net313),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[16][1] ));
 DLH_X1 _11782_ (.D(net304),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[16][2] ));
 DLH_X1 _11783_ (.D(net299),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[16][3] ));
 DLH_X1 _11784_ (.D(net294),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[16][4] ));
 DLH_X1 _11785_ (.D(net288),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[16][5] ));
 DLH_X1 _11786_ (.D(net282),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[16][6] ));
 DLH_X1 _11787_ (.D(net276),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[16][7] ));
 DLH_X1 _11788_ (.D(net316),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[24][0] ));
 DLH_X1 _11789_ (.D(net313),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[24][1] ));
 DLH_X1 _11790_ (.D(net304),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[24][2] ));
 DLH_X1 _11791_ (.D(net299),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[24][3] ));
 DLH_X1 _11792_ (.D(net294),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[24][4] ));
 DLH_X1 _11793_ (.D(net288),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[24][5] ));
 DLH_X1 _11794_ (.D(net282),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[24][6] ));
 DLH_X1 _11795_ (.D(net276),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[24][7] ));
 DLH_X1 _11796_ (.D(net316),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[4][0] ));
 DLH_X1 _11797_ (.D(net312),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[4][1] ));
 DLH_X1 _11798_ (.D(net304),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[4][2] ));
 DLH_X1 _11799_ (.D(net299),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[4][3] ));
 DLH_X1 _11800_ (.D(net294),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[4][4] ));
 DLH_X1 _11801_ (.D(net288),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[4][5] ));
 DLH_X1 _11802_ (.D(net282),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[4][6] ));
 DLH_X1 _11803_ (.D(net276),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[4][7] ));
 DLH_X1 _11804_ (.D(net316),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[15][0] ));
 DLH_X1 _11805_ (.D(net313),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[15][1] ));
 DLH_X1 _11806_ (.D(net304),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[15][2] ));
 DLH_X1 _11807_ (.D(net299),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[15][3] ));
 DLH_X1 _11808_ (.D(net294),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[15][4] ));
 DLH_X1 _11809_ (.D(net288),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[15][5] ));
 DLH_X1 _11810_ (.D(net282),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[15][6] ));
 DLH_X1 _11811_ (.D(net276),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[15][7] ));
 DLH_X1 _11812_ (.D(net316),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[11][0] ));
 DLH_X1 _11813_ (.D(net312),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[11][1] ));
 DLH_X1 _11814_ (.D(net304),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[11][2] ));
 DLH_X1 _11815_ (.D(net298),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[11][3] ));
 DLH_X1 _11816_ (.D(net294),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[11][4] ));
 DLH_X1 _11817_ (.D(net288),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[11][5] ));
 DLH_X1 _11818_ (.D(net282),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[11][6] ));
 DLH_X1 _11819_ (.D(net276),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[11][7] ));
 DLH_X1 _11820_ (.D(net316),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[5][0] ));
 DLH_X1 _11821_ (.D(net312),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[5][1] ));
 DLH_X1 _11822_ (.D(net304),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[5][2] ));
 DLH_X1 _11823_ (.D(net299),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[5][3] ));
 DLH_X1 _11824_ (.D(net294),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[5][4] ));
 DLH_X1 _11825_ (.D(net288),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[5][5] ));
 DLH_X1 _11826_ (.D(net282),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[5][6] ));
 DLH_X1 _11827_ (.D(net276),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[5][7] ));
 DLH_X1 _11828_ (.D(net316),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[23][0] ));
 DLH_X1 _11829_ (.D(net312),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[23][1] ));
 DLH_X1 _11830_ (.D(net304),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[23][2] ));
 DLH_X1 _11831_ (.D(net299),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[23][3] ));
 DLH_X1 _11832_ (.D(net294),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[23][4] ));
 DLH_X1 _11833_ (.D(net288),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[23][5] ));
 DLH_X1 _11834_ (.D(net282),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[23][6] ));
 DLH_X1 _11835_ (.D(net276),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[23][7] ));
 DLH_X1 _11836_ (.D(net316),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[19][0] ));
 DLH_X1 _11837_ (.D(net313),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[19][1] ));
 DLH_X1 _11838_ (.D(net304),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[19][2] ));
 DLH_X1 _11839_ (.D(net299),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[19][3] ));
 DLH_X1 _11840_ (.D(net294),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[19][4] ));
 DLH_X1 _11841_ (.D(net288),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[19][5] ));
 DLH_X1 _11842_ (.D(net282),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[19][6] ));
 DLH_X1 _11843_ (.D(net276),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[19][7] ));
 DLH_X1 _11844_ (.D(net316),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[31][0] ));
 DLH_X1 _11845_ (.D(net313),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[31][1] ));
 DLH_X1 _11846_ (.D(net304),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[31][2] ));
 DLH_X1 _11847_ (.D(net298),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[31][3] ));
 DLH_X1 _11848_ (.D(net294),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[31][4] ));
 DLH_X1 _11849_ (.D(net288),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[31][5] ));
 DLH_X1 _11850_ (.D(net282),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[31][6] ));
 DLH_X1 _11851_ (.D(net276),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[31][7] ));
 DLH_X1 _11852_ (.D(net316),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[6][0] ));
 DLH_X1 _11853_ (.D(net312),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[6][1] ));
 DLH_X1 _11854_ (.D(net304),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[6][2] ));
 DLH_X1 _11855_ (.D(net299),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[6][3] ));
 DLH_X1 _11856_ (.D(net294),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[6][4] ));
 DLH_X1 _11857_ (.D(net288),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[6][5] ));
 DLH_X1 _11858_ (.D(net282),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[6][6] ));
 DLH_X1 _11859_ (.D(net276),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[6][7] ));
 DLH_X1 _11860_ (.D(net316),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[14][0] ));
 DLH_X1 _11861_ (.D(net313),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[14][1] ));
 DLH_X1 _11862_ (.D(net304),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[14][2] ));
 DLH_X1 _11863_ (.D(net299),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[14][3] ));
 DLH_X1 _11864_ (.D(net294),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[14][4] ));
 DLH_X1 _11865_ (.D(net288),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[14][5] ));
 DLH_X1 _11866_ (.D(net282),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[14][6] ));
 DLH_X1 _11867_ (.D(net276),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[14][7] ));
 DLH_X1 _11868_ (.D(net316),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[30][0] ));
 DLH_X1 _11869_ (.D(net312),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[30][1] ));
 DLH_X1 _11870_ (.D(net304),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[30][2] ));
 DLH_X1 _11871_ (.D(net298),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[30][3] ));
 DLH_X1 _11872_ (.D(net294),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[30][4] ));
 DLH_X1 _11873_ (.D(net288),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[30][5] ));
 DLH_X1 _11874_ (.D(net282),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[30][6] ));
 DLH_X1 _11875_ (.D(net276),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[30][7] ));
 DLH_X1 _11876_ (.D(net316),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[22][0] ));
 DLH_X1 _11877_ (.D(net313),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[22][1] ));
 DLH_X1 _11878_ (.D(net305),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[22][2] ));
 DLH_X1 _11879_ (.D(net299),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[22][3] ));
 DLH_X1 _11880_ (.D(net294),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[22][4] ));
 DLH_X1 _11881_ (.D(net288),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[22][5] ));
 DLH_X1 _11882_ (.D(net282),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[22][6] ));
 DLH_X1 _11883_ (.D(net276),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[22][7] ));
 DLH_X1 _11884_ (.D(net316),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[7][0] ));
 DLH_X1 _11885_ (.D(net313),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[7][1] ));
 DLH_X1 _11886_ (.D(net304),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[7][2] ));
 DLH_X1 _11887_ (.D(net298),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[7][3] ));
 DLH_X1 _11888_ (.D(net294),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[7][4] ));
 DLH_X1 _11889_ (.D(net288),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[7][5] ));
 DLH_X1 _11890_ (.D(net282),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[7][6] ));
 DLH_X1 _11891_ (.D(net276),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[7][7] ));
 DLH_X1 _11892_ (.D(net316),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[29][0] ));
 DLH_X1 _11893_ (.D(net312),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[29][1] ));
 DLH_X1 _11894_ (.D(net304),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[29][2] ));
 DLH_X1 _11895_ (.D(net299),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[29][3] ));
 DLH_X1 _11896_ (.D(net294),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[29][4] ));
 DLH_X1 _11897_ (.D(net288),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[29][5] ));
 DLH_X1 _11898_ (.D(net282),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[29][6] ));
 DLH_X1 _11899_ (.D(net276),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[29][7] ));
 DLH_X1 _11900_ (.D(net316),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[12][0] ));
 DLH_X1 _11901_ (.D(net312),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[12][1] ));
 DLH_X1 _11902_ (.D(net304),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[12][2] ));
 DLH_X1 _11903_ (.D(net299),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[12][3] ));
 DLH_X1 _11904_ (.D(net294),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[12][4] ));
 DLH_X1 _11905_ (.D(net288),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[12][5] ));
 DLH_X1 _11906_ (.D(net282),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[12][6] ));
 DLH_X1 _11907_ (.D(net276),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[12][7] ));
 DLH_X1 _11908_ (.D(net316),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[17][0] ));
 DLH_X1 _11909_ (.D(net313),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[17][1] ));
 DLH_X1 _11910_ (.D(net305),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[17][2] ));
 DLH_X1 _11911_ (.D(net298),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[17][3] ));
 DLH_X1 _11912_ (.D(net294),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[17][4] ));
 DLH_X1 _11913_ (.D(net288),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[17][5] ));
 DLH_X1 _11914_ (.D(net282),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[17][6] ));
 DLH_X1 _11915_ (.D(net276),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[17][7] ));
 DLH_X1 _11916_ (.D(net316),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[28][0] ));
 DLH_X1 _11917_ (.D(net312),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[28][1] ));
 DLH_X1 _11918_ (.D(net304),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[28][2] ));
 DLH_X1 _11919_ (.D(net299),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[28][3] ));
 DLH_X1 _11920_ (.D(net294),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[28][4] ));
 DLH_X1 _11921_ (.D(net288),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[28][5] ));
 DLH_X1 _11922_ (.D(net282),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[28][6] ));
 DLH_X1 _11923_ (.D(net276),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[28][7] ));
 DLH_X1 _11924_ (.D(net316),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[8][0] ));
 DLH_X1 _11925_ (.D(net312),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[8][1] ));
 DLH_X1 _11926_ (.D(net304),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[8][2] ));
 DLH_X1 _11927_ (.D(net299),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[8][3] ));
 DLH_X1 _11928_ (.D(net294),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[8][4] ));
 DLH_X1 _11929_ (.D(net288),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[8][5] ));
 DLH_X1 _11930_ (.D(net282),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[8][6] ));
 DLH_X1 _11931_ (.D(net276),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[8][7] ));
 DLH_X1 _11932_ (.D(net316),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[21][0] ));
 DLH_X1 _11933_ (.D(net313),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[21][1] ));
 DLH_X1 _11934_ (.D(net304),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[21][2] ));
 DLH_X1 _11935_ (.D(net299),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[21][3] ));
 DLH_X1 _11936_ (.D(net294),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[21][4] ));
 DLH_X1 _11937_ (.D(net288),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[21][5] ));
 DLH_X1 _11938_ (.D(net282),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[21][6] ));
 DLH_X1 _11939_ (.D(net276),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[21][7] ));
 DLH_X1 _11940_ (.D(net316),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[27][0] ));
 DLH_X1 _11941_ (.D(net312),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[27][1] ));
 DLH_X1 _11942_ (.D(net305),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[27][2] ));
 DLH_X1 _11943_ (.D(net298),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[27][3] ));
 DLH_X1 _11944_ (.D(net294),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[27][4] ));
 DLH_X1 _11945_ (.D(net288),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[27][5] ));
 DLH_X1 _11946_ (.D(net282),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[27][6] ));
 DLH_X1 _11947_ (.D(net276),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[27][7] ));
 DLH_X1 _11948_ (.D(net316),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[18][0] ));
 DLH_X1 _11949_ (.D(net313),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[18][1] ));
 DLH_X1 _11950_ (.D(net305),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[18][2] ));
 DLH_X1 _11951_ (.D(net299),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[18][3] ));
 DLH_X1 _11952_ (.D(net294),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[18][4] ));
 DLH_X1 _11953_ (.D(net288),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[18][5] ));
 DLH_X1 _11954_ (.D(net282),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[18][6] ));
 DLH_X1 _11955_ (.D(net276),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.mem[18][7] ));
 DLL_X1 _11956_ (.D(\lut.gen_sub_units_scm.__8.sub_unit_i.cg_we_global.en_i ),
    .GN(clknet_level_5_1_114__00532_),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.cg_we_global.clk_en ));
 DLL_X1 _11957_ (.D(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__0.cg_i.en_i ),
    .GN(clknet_level_2_1_862__00555_),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_en ));
 DLL_X1 _11958_ (.D(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__1.cg_i.en_i ),
    .GN(clknet_level_2_1_141__00555_),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_en ));
 DLL_X1 _11959_ (.D(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__2.cg_i.en_i ),
    .GN(clknet_level_2_1_450__00555_),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_en ));
 DLL_X1 _11960_ (.D(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__3.cg_i.en_i ),
    .GN(clknet_level_2_1_862__00555_),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_en ));
 DLL_X1 _11961_ (.D(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__4.cg_i.en_i ),
    .GN(clknet_level_2_1_244__00555_),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_en ));
 DLL_X1 _11962_ (.D(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__5.cg_i.en_i ),
    .GN(clknet_level_2_1_244__00555_),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_en ));
 DLL_X1 _11963_ (.D(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__6.cg_i.en_i ),
    .GN(clknet_level_2_1_553__00555_),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_en ));
 DLL_X1 _11964_ (.D(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__7.cg_i.en_i ),
    .GN(clknet_level_2_1_450__00555_),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_en ));
 DLL_X1 _11965_ (.D(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__8.cg_i.en_i ),
    .GN(clknet_level_2_1_244__00555_),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_en ));
 DLL_X1 _11966_ (.D(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__9.cg_i.en_i ),
    .GN(clknet_level_2_1_656__00555_),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_en ));
 DLL_X1 _11967_ (.D(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__10.cg_i.en_i ),
    .GN(clknet_level_2_1_656__00555_),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_en ));
 DLL_X1 _11968_ (.D(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__11.cg_i.en_i ),
    .GN(clknet_level_2_1_759__00555_),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_en ));
 DLL_X1 _11969_ (.D(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__12.cg_i.en_i ),
    .GN(clknet_level_2_1_450__00555_),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_en ));
 DLL_X1 _11970_ (.D(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__13.cg_i.en_i ),
    .GN(clknet_level_2_1_141__00555_),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_en ));
 DLL_X1 _11971_ (.D(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__14.cg_i.en_i ),
    .GN(clknet_level_2_1_347__00555_),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_en ));
 DLL_X1 _11972_ (.D(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__15.cg_i.en_i ),
    .GN(clknet_level_2_1_347__00555_),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_en ));
 DLL_X1 _11973_ (.D(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__16.cg_i.en_i ),
    .GN(clknet_level_2_1_347__00555_),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_en ));
 DLL_X1 _11974_ (.D(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__17.cg_i.en_i ),
    .GN(clknet_level_2_1_759__00555_),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_en ));
 DLL_X1 _11975_ (.D(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__18.cg_i.en_i ),
    .GN(clknet_level_2_1_347__00555_),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_en ));
 DLL_X1 _11976_ (.D(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__19.cg_i.en_i ),
    .GN(clknet_level_2_1_141__00555_),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_en ));
 DLL_X1 _11977_ (.D(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__20.cg_i.en_i ),
    .GN(clknet_level_2_1_141__00555_),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_en ));
 DLL_X1 _11978_ (.D(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__21.cg_i.en_i ),
    .GN(clknet_level_2_1_862__00555_),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_en ));
 DLL_X1 _11979_ (.D(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__22.cg_i.en_i ),
    .GN(clknet_level_2_1_347__00555_),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_en ));
 DLL_X1 _11980_ (.D(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__23.cg_i.en_i ),
    .GN(clknet_level_2_1_244__00555_),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_en ));
 DLL_X1 _11981_ (.D(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__24.cg_i.en_i ),
    .GN(clknet_level_2_1_450__00555_),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_en ));
 DLL_X1 _11982_ (.D(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__25.cg_i.en_i ),
    .GN(clknet_level_2_1_656__00555_),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_en ));
 DLL_X1 _11983_ (.D(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__26.cg_i.en_i ),
    .GN(clknet_level_2_1_141__00555_),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_en ));
 DLL_X1 _11984_ (.D(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__27.cg_i.en_i ),
    .GN(clknet_level_2_1_759__00555_),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_en ));
 DLL_X1 _11985_ (.D(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__28.cg_i.en_i ),
    .GN(clknet_level_2_1_656__00555_),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_en ));
 DLL_X1 _11986_ (.D(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__29.cg_i.en_i ),
    .GN(clknet_level_2_1_450__00555_),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_en ));
 DLL_X1 _11987_ (.D(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__30.cg_i.en_i ),
    .GN(clknet_level_2_1_553__00555_),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_en ));
 DLL_X1 _11988_ (.D(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__31.cg_i.en_i ),
    .GN(clknet_level_2_1_553__00555_),
    .Q(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_en ));
 DLH_X1 _11989_ (.D(net319),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[13][0] ));
 DLH_X1 _11990_ (.D(net314),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[13][1] ));
 DLH_X1 _11991_ (.D(net309),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[13][2] ));
 DLH_X1 _11992_ (.D(net301),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[13][3] ));
 DLH_X1 _11993_ (.D(net296),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[13][4] ));
 DLH_X1 _11994_ (.D(net290),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[13][5] ));
 DLH_X1 _11995_ (.D(net286),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[13][6] ));
 DLH_X1 _11996_ (.D(net278),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[13][7] ));
 DLH_X1 _11997_ (.D(net318),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[1][0] ));
 DLH_X1 _11998_ (.D(net314),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[1][1] ));
 DLH_X1 _11999_ (.D(net309),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[1][2] ));
 DLH_X1 _12000_ (.D(net301),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[1][3] ));
 DLH_X1 _12001_ (.D(net296),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[1][4] ));
 DLH_X1 _12002_ (.D(net290),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[1][5] ));
 DLH_X1 _12003_ (.D(net286),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[1][6] ));
 DLH_X1 _12004_ (.D(net278),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[1][7] ));
 DLH_X1 _12005_ (.D(net318),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[26][0] ));
 DLH_X1 _12006_ (.D(net314),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[26][1] ));
 DLH_X1 _12007_ (.D(net309),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[26][2] ));
 DLH_X1 _12008_ (.D(net301),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[26][3] ));
 DLH_X1 _12009_ (.D(net296),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[26][4] ));
 DLH_X1 _12010_ (.D(net289),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[26][5] ));
 DLH_X1 _12011_ (.D(net286),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[26][6] ));
 DLH_X1 _12012_ (.D(net278),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[26][7] ));
 DLH_X1 _12013_ (.D(net318),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[9][0] ));
 DLH_X1 _12014_ (.D(net314),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[9][1] ));
 DLH_X1 _12015_ (.D(net309),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[9][2] ));
 DLH_X1 _12016_ (.D(net301),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[9][3] ));
 DLH_X1 _12017_ (.D(net296),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[9][4] ));
 DLH_X1 _12018_ (.D(net289),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[9][5] ));
 DLH_X1 _12019_ (.D(net286),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[9][6] ));
 DLH_X1 _12020_ (.D(net278),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[9][7] ));
 DLH_X1 _12021_ (.D(net319),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[0][0] ));
 DLH_X1 _12022_ (.D(net312),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[0][1] ));
 DLH_X1 _12023_ (.D(net304),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[0][2] ));
 DLH_X1 _12024_ (.D(net303),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[0][3] ));
 DLH_X1 _12025_ (.D(net295),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[0][4] ));
 DLH_X1 _12026_ (.D(net292),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[0][5] ));
 DLH_X1 _12027_ (.D(net285),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[0][6] ));
 DLH_X1 _12028_ (.D(net279),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[0][7] ));
 DLH_X1 _12029_ (.D(net319),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[20][0] ));
 DLH_X1 _12030_ (.D(net314),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[20][1] ));
 DLH_X1 _12031_ (.D(net309),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[20][2] ));
 DLH_X1 _12032_ (.D(net301),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[20][3] ));
 DLH_X1 _12033_ (.D(net296),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[20][4] ));
 DLH_X1 _12034_ (.D(net289),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[20][5] ));
 DLH_X1 _12035_ (.D(net286),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[20][6] ));
 DLH_X1 _12036_ (.D(net278),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[20][7] ));
 DLH_X1 _12037_ (.D(net318),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[2][0] ));
 DLH_X1 _12038_ (.D(net314),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[2][1] ));
 DLH_X1 _12039_ (.D(net307),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[2][2] ));
 DLH_X1 _12040_ (.D(net301),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[2][3] ));
 DLH_X1 _12041_ (.D(net296),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[2][4] ));
 DLH_X1 _12042_ (.D(net289),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[2][5] ));
 DLH_X1 _12043_ (.D(net281),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[2][6] ));
 DLH_X1 _12044_ (.D(net278),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[2][7] ));
 DLH_X1 _12045_ (.D(net319),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[25][0] ));
 DLH_X1 _12046_ (.D(net312),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[25][1] ));
 DLH_X1 _12047_ (.D(net309),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[25][2] ));
 DLH_X1 _12048_ (.D(net301),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[25][3] ));
 DLH_X1 _12049_ (.D(net296),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[25][4] ));
 DLH_X1 _12050_ (.D(net290),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[25][5] ));
 DLH_X1 _12051_ (.D(net286),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[25][6] ));
 DLH_X1 _12052_ (.D(net278),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[25][7] ));
 DLH_X1 _12053_ (.D(net318),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[10][0] ));
 DLH_X1 _12054_ (.D(net314),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[10][1] ));
 DLH_X1 _12055_ (.D(net307),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[10][2] ));
 DLH_X1 _12056_ (.D(net301),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[10][3] ));
 DLH_X1 _12057_ (.D(net296),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[10][4] ));
 DLH_X1 _12058_ (.D(net289),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[10][5] ));
 DLH_X1 _12059_ (.D(net286),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[10][6] ));
 DLH_X1 _12060_ (.D(net278),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[10][7] ));
 DLH_X1 _12061_ (.D(net318),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[3][0] ));
 DLH_X1 _12062_ (.D(net314),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[3][1] ));
 DLH_X1 _12063_ (.D(net309),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[3][2] ));
 DLH_X1 _12064_ (.D(net301),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[3][3] ));
 DLH_X1 _12065_ (.D(net296),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[3][4] ));
 DLH_X1 _12066_ (.D(net289),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[3][5] ));
 DLH_X1 _12067_ (.D(net281),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[3][6] ));
 DLH_X1 _12068_ (.D(net278),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[3][7] ));
 DLH_X1 _12069_ (.D(net318),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[16][0] ));
 DLH_X1 _12070_ (.D(net314),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[16][1] ));
 DLH_X1 _12071_ (.D(net307),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[16][2] ));
 DLH_X1 _12072_ (.D(net301),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[16][3] ));
 DLH_X1 _12073_ (.D(net296),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[16][4] ));
 DLH_X1 _12074_ (.D(net289),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[16][5] ));
 DLH_X1 _12075_ (.D(net286),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[16][6] ));
 DLH_X1 _12076_ (.D(net278),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[16][7] ));
 DLH_X1 _12077_ (.D(net318),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[24][0] ));
 DLH_X1 _12078_ (.D(net314),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[24][1] ));
 DLH_X1 _12079_ (.D(net307),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[24][2] ));
 DLH_X1 _12080_ (.D(net301),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[24][3] ));
 DLH_X1 _12081_ (.D(net296),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[24][4] ));
 DLH_X1 _12082_ (.D(net290),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[24][5] ));
 DLH_X1 _12083_ (.D(net281),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[24][6] ));
 DLH_X1 _12084_ (.D(net278),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[24][7] ));
 DLH_X1 _12085_ (.D(net319),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[4][0] ));
 DLH_X1 _12086_ (.D(net314),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[4][1] ));
 DLH_X1 _12087_ (.D(net307),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[4][2] ));
 DLH_X1 _12088_ (.D(net301),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[4][3] ));
 DLH_X1 _12089_ (.D(net296),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[4][4] ));
 DLH_X1 _12090_ (.D(net289),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[4][5] ));
 DLH_X1 _12091_ (.D(net281),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[4][6] ));
 DLH_X1 _12092_ (.D(net278),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[4][7] ));
 DLH_X1 _12093_ (.D(net318),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[15][0] ));
 DLH_X1 _12094_ (.D(net314),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[15][1] ));
 DLH_X1 _12095_ (.D(net309),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[15][2] ));
 DLH_X1 _12096_ (.D(net301),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[15][3] ));
 DLH_X1 _12097_ (.D(net296),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[15][4] ));
 DLH_X1 _12098_ (.D(net289),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[15][5] ));
 DLH_X1 _12099_ (.D(net286),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[15][6] ));
 DLH_X1 _12100_ (.D(net278),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[15][7] ));
 DLH_X1 _12101_ (.D(net318),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[11][0] ));
 DLH_X1 _12102_ (.D(net314),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[11][1] ));
 DLH_X1 _12103_ (.D(net307),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[11][2] ));
 DLH_X1 _12104_ (.D(net301),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[11][3] ));
 DLH_X1 _12105_ (.D(net296),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[11][4] ));
 DLH_X1 _12106_ (.D(net289),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[11][5] ));
 DLH_X1 _12107_ (.D(net286),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[11][6] ));
 DLH_X1 _12108_ (.D(net278),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[11][7] ));
 DLH_X1 _12109_ (.D(net318),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[5][0] ));
 DLH_X1 _12110_ (.D(net314),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[5][1] ));
 DLH_X1 _12111_ (.D(net307),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[5][2] ));
 DLH_X1 _12112_ (.D(net301),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[5][3] ));
 DLH_X1 _12113_ (.D(net296),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[5][4] ));
 DLH_X1 _12114_ (.D(net290),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[5][5] ));
 DLH_X1 _12115_ (.D(net286),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[5][6] ));
 DLH_X1 _12116_ (.D(net278),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[5][7] ));
 DLH_X1 _12117_ (.D(net319),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[23][0] ));
 DLH_X1 _12118_ (.D(net314),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[23][1] ));
 DLH_X1 _12119_ (.D(net309),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[23][2] ));
 DLH_X1 _12120_ (.D(net301),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[23][3] ));
 DLH_X1 _12121_ (.D(net296),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[23][4] ));
 DLH_X1 _12122_ (.D(net290),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[23][5] ));
 DLH_X1 _12123_ (.D(net286),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[23][6] ));
 DLH_X1 _12124_ (.D(net278),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[23][7] ));
 DLH_X1 _12125_ (.D(net318),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[19][0] ));
 DLH_X1 _12126_ (.D(net314),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[19][1] ));
 DLH_X1 _12127_ (.D(net309),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[19][2] ));
 DLH_X1 _12128_ (.D(net301),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[19][3] ));
 DLH_X1 _12129_ (.D(net296),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[19][4] ));
 DLH_X1 _12130_ (.D(net289),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[19][5] ));
 DLH_X1 _12131_ (.D(net281),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[19][6] ));
 DLH_X1 _12132_ (.D(net278),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[19][7] ));
 DLH_X1 _12133_ (.D(net318),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[31][0] ));
 DLH_X1 _12134_ (.D(net314),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[31][1] ));
 DLH_X1 _12135_ (.D(net307),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[31][2] ));
 DLH_X1 _12136_ (.D(net301),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[31][3] ));
 DLH_X1 _12137_ (.D(net296),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[31][4] ));
 DLH_X1 _12138_ (.D(net289),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[31][5] ));
 DLH_X1 _12139_ (.D(net286),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[31][6] ));
 DLH_X1 _12140_ (.D(net278),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[31][7] ));
 DLH_X1 _12141_ (.D(net318),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[6][0] ));
 DLH_X1 _12142_ (.D(net314),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[6][1] ));
 DLH_X1 _12143_ (.D(net309),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[6][2] ));
 DLH_X1 _12144_ (.D(net301),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[6][3] ));
 DLH_X1 _12145_ (.D(net296),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[6][4] ));
 DLH_X1 _12146_ (.D(net289),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[6][5] ));
 DLH_X1 _12147_ (.D(net286),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[6][6] ));
 DLH_X1 _12148_ (.D(net278),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[6][7] ));
 DLH_X1 _12149_ (.D(net318),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[14][0] ));
 DLH_X1 _12150_ (.D(net314),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[14][1] ));
 DLH_X1 _12151_ (.D(net309),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[14][2] ));
 DLH_X1 _12152_ (.D(net301),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[14][3] ));
 DLH_X1 _12153_ (.D(net296),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[14][4] ));
 DLH_X1 _12154_ (.D(net289),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[14][5] ));
 DLH_X1 _12155_ (.D(net286),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[14][6] ));
 DLH_X1 _12156_ (.D(net278),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[14][7] ));
 DLH_X1 _12157_ (.D(net318),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[30][0] ));
 DLH_X1 _12158_ (.D(net314),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[30][1] ));
 DLH_X1 _12159_ (.D(net304),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[30][2] ));
 DLH_X1 _12160_ (.D(net301),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[30][3] ));
 DLH_X1 _12161_ (.D(net296),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[30][4] ));
 DLH_X1 _12162_ (.D(net289),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[30][5] ));
 DLH_X1 _12163_ (.D(net286),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[30][6] ));
 DLH_X1 _12164_ (.D(net278),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[30][7] ));
 DLH_X1 _12165_ (.D(net318),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[22][0] ));
 DLH_X1 _12166_ (.D(net312),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[22][1] ));
 DLH_X1 _12167_ (.D(net307),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[22][2] ));
 DLH_X1 _12168_ (.D(net301),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[22][3] ));
 DLH_X1 _12169_ (.D(net296),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[22][4] ));
 DLH_X1 _12170_ (.D(net289),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[22][5] ));
 DLH_X1 _12171_ (.D(net281),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[22][6] ));
 DLH_X1 _12172_ (.D(net278),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[22][7] ));
 DLH_X1 _12173_ (.D(net319),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[7][0] ));
 DLH_X1 _12174_ (.D(net314),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[7][1] ));
 DLH_X1 _12175_ (.D(net307),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[7][2] ));
 DLH_X1 _12176_ (.D(net301),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[7][3] ));
 DLH_X1 _12177_ (.D(net296),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[7][4] ));
 DLH_X1 _12178_ (.D(net289),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[7][5] ));
 DLH_X1 _12179_ (.D(net286),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[7][6] ));
 DLH_X1 _12180_ (.D(net278),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[7][7] ));
 DLH_X1 _12181_ (.D(net318),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[29][0] ));
 DLH_X1 _12182_ (.D(net314),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[29][1] ));
 DLH_X1 _12183_ (.D(net309),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[29][2] ));
 DLH_X1 _12184_ (.D(net301),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[29][3] ));
 DLH_X1 _12185_ (.D(net296),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[29][4] ));
 DLH_X1 _12186_ (.D(net290),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[29][5] ));
 DLH_X1 _12187_ (.D(net286),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[29][6] ));
 DLH_X1 _12188_ (.D(net278),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[29][7] ));
 DLH_X1 _12189_ (.D(net318),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[12][0] ));
 DLH_X1 _12190_ (.D(net314),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[12][1] ));
 DLH_X1 _12191_ (.D(net307),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[12][2] ));
 DLH_X1 _12192_ (.D(net301),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[12][3] ));
 DLH_X1 _12193_ (.D(net296),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[12][4] ));
 DLH_X1 _12194_ (.D(net289),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[12][5] ));
 DLH_X1 _12195_ (.D(net286),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[12][6] ));
 DLH_X1 _12196_ (.D(net278),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[12][7] ));
 DLH_X1 _12197_ (.D(net318),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[17][0] ));
 DLH_X1 _12198_ (.D(net314),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[17][1] ));
 DLH_X1 _12199_ (.D(net304),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[17][2] ));
 DLH_X1 _12200_ (.D(net301),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[17][3] ));
 DLH_X1 _12201_ (.D(net296),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[17][4] ));
 DLH_X1 _12202_ (.D(net289),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[17][5] ));
 DLH_X1 _12203_ (.D(net281),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[17][6] ));
 DLH_X1 _12204_ (.D(net278),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[17][7] ));
 DLH_X1 _12205_ (.D(net318),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[28][0] ));
 DLH_X1 _12206_ (.D(net314),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[28][1] ));
 DLH_X1 _12207_ (.D(net307),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[28][2] ));
 DLH_X1 _12208_ (.D(net301),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[28][3] ));
 DLH_X1 _12209_ (.D(net296),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[28][4] ));
 DLH_X1 _12210_ (.D(net289),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[28][5] ));
 DLH_X1 _12211_ (.D(net286),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[28][6] ));
 DLH_X1 _12212_ (.D(net278),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[28][7] ));
 DLH_X1 _12213_ (.D(net318),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[8][0] ));
 DLH_X1 _12214_ (.D(net314),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[8][1] ));
 DLH_X1 _12215_ (.D(net309),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[8][2] ));
 DLH_X1 _12216_ (.D(net301),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[8][3] ));
 DLH_X1 _12217_ (.D(net296),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[8][4] ));
 DLH_X1 _12218_ (.D(net289),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[8][5] ));
 DLH_X1 _12219_ (.D(net281),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[8][6] ));
 DLH_X1 _12220_ (.D(net278),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[8][7] ));
 DLH_X1 _12221_ (.D(net318),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[21][0] ));
 DLH_X1 _12222_ (.D(net314),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[21][1] ));
 DLH_X1 _12223_ (.D(net307),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[21][2] ));
 DLH_X1 _12224_ (.D(net301),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[21][3] ));
 DLH_X1 _12225_ (.D(net296),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[21][4] ));
 DLH_X1 _12226_ (.D(net290),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[21][5] ));
 DLH_X1 _12227_ (.D(net281),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[21][6] ));
 DLH_X1 _12228_ (.D(net278),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[21][7] ));
 DLH_X1 _12229_ (.D(net319),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[27][0] ));
 DLH_X1 _12230_ (.D(net314),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[27][1] ));
 DLH_X1 _12231_ (.D(net309),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[27][2] ));
 DLH_X1 _12232_ (.D(net301),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[27][3] ));
 DLH_X1 _12233_ (.D(net296),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[27][4] ));
 DLH_X1 _12234_ (.D(net289),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[27][5] ));
 DLH_X1 _12235_ (.D(net286),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[27][6] ));
 DLH_X1 _12236_ (.D(net278),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[27][7] ));
 DLH_X1 _12237_ (.D(net319),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[18][0] ));
 DLH_X1 _12238_ (.D(net314),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[18][1] ));
 DLH_X1 _12239_ (.D(net309),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[18][2] ));
 DLH_X1 _12240_ (.D(net301),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[18][3] ));
 DLH_X1 _12241_ (.D(net296),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[18][4] ));
 DLH_X1 _12242_ (.D(net289),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[18][5] ));
 DLH_X1 _12243_ (.D(net286),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[18][6] ));
 DLH_X1 _12244_ (.D(net278),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.mem[18][7] ));
 DLL_X1 _12245_ (.D(\lut.gen_sub_units_scm.__7.sub_unit_i.cg_we_global.en_i ),
    .GN(clknet_level_5_1_2116__00532_),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.cg_we_global.clk_en ));
 DLL_X1 _12246_ (.D(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__0.cg_i.en_i ),
    .GN(clknet_level_2_1_680__00558_),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_en ));
 DLL_X1 _12247_ (.D(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__1.cg_i.en_i ),
    .GN(clknet_level_2_1_474__00558_),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_en ));
 DLL_X1 _12248_ (.D(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__2.cg_i.en_i ),
    .GN(clknet_level_2_1_165__00558_),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_en ));
 DLL_X1 _12249_ (.D(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__3.cg_i.en_i ),
    .GN(clknet_level_2_1_886__00558_),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_en ));
 DLL_X1 _12250_ (.D(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__4.cg_i.en_i ),
    .GN(clknet_level_2_1_268__00558_),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_en ));
 DLL_X1 _12251_ (.D(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__5.cg_i.en_i ),
    .GN(clknet_level_2_1_680__00558_),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_en ));
 DLL_X1 _12252_ (.D(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__6.cg_i.en_i ),
    .GN(clknet_level_2_1_783__00558_),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_en ));
 DLL_X1 _12253_ (.D(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__7.cg_i.en_i ),
    .GN(clknet_level_2_1_268__00558_),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_en ));
 DLL_X1 _12254_ (.D(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__8.cg_i.en_i ),
    .GN(clknet_level_2_1_371__00558_),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_en ));
 DLL_X1 _12255_ (.D(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__9.cg_i.en_i ),
    .GN(clknet_level_2_1_886__00558_),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_en ));
 DLL_X1 _12256_ (.D(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__10.cg_i.en_i ),
    .GN(clknet_level_2_1_680__00558_),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_en ));
 DLL_X1 _12257_ (.D(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__11.cg_i.en_i ),
    .GN(clknet_level_2_1_577__00558_),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_en ));
 DLL_X1 _12258_ (.D(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__12.cg_i.en_i ),
    .GN(clknet_level_2_1_268__00558_),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_en ));
 DLL_X1 _12259_ (.D(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__13.cg_i.en_i ),
    .GN(clknet_level_2_1_886__00558_),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_en ));
 DLL_X1 _12260_ (.D(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__14.cg_i.en_i ),
    .GN(clknet_level_2_1_474__00558_),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_en ));
 DLL_X1 _12261_ (.D(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__15.cg_i.en_i ),
    .GN(clknet_level_2_1_783__00558_),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_en ));
 DLL_X1 _12262_ (.D(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__16.cg_i.en_i ),
    .GN(clknet_level_2_1_680__00558_),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_en ));
 DLL_X1 _12263_ (.D(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__17.cg_i.en_i ),
    .GN(clknet_level_2_1_577__00558_),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_en ));
 DLL_X1 _12264_ (.D(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__18.cg_i.en_i ),
    .GN(clknet_level_2_1_474__00558_),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_en ));
 DLL_X1 _12265_ (.D(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__19.cg_i.en_i ),
    .GN(clknet_level_2_1_474__00558_),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_en ));
 DLL_X1 _12266_ (.D(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__20.cg_i.en_i ),
    .GN(clknet_level_2_1_474__00558_),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_en ));
 DLL_X1 _12267_ (.D(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__21.cg_i.en_i ),
    .GN(clknet_level_2_1_680__00558_),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_en ));
 DLL_X1 _12268_ (.D(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__22.cg_i.en_i ),
    .GN(clknet_level_2_1_577__00558_),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_en ));
 DLL_X1 _12269_ (.D(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__23.cg_i.en_i ),
    .GN(clknet_level_2_1_371__00558_),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_en ));
 DLL_X1 _12270_ (.D(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__24.cg_i.en_i ),
    .GN(clknet_level_2_1_268__00558_),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_en ));
 DLL_X1 _12271_ (.D(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__25.cg_i.en_i ),
    .GN(clknet_level_2_1_680__00558_),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_en ));
 DLL_X1 _12272_ (.D(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__26.cg_i.en_i ),
    .GN(clknet_level_2_1_371__00558_),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_en ));
 DLL_X1 _12273_ (.D(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__27.cg_i.en_i ),
    .GN(clknet_level_2_1_371__00558_),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_en ));
 DLL_X1 _12274_ (.D(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__28.cg_i.en_i ),
    .GN(clknet_level_2_1_886__00558_),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_en ));
 DLL_X1 _12275_ (.D(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__29.cg_i.en_i ),
    .GN(clknet_level_2_1_886__00558_),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_en ));
 DLL_X1 _12276_ (.D(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__30.cg_i.en_i ),
    .GN(clknet_level_2_1_268__00558_),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_en ));
 DLL_X1 _12277_ (.D(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__31.cg_i.en_i ),
    .GN(clknet_level_2_1_680__00558_),
    .Q(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_en ));
 DLH_X1 _12278_ (.D(net316),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[13][0] ));
 DLH_X1 _12279_ (.D(net312),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[13][1] ));
 DLH_X1 _12280_ (.D(net304),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[13][2] ));
 DLH_X1 _12281_ (.D(net298),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[13][3] ));
 DLH_X1 _12282_ (.D(net295),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[13][4] ));
 DLH_X1 _12283_ (.D(net288),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[13][5] ));
 DLH_X1 _12284_ (.D(net282),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[13][6] ));
 DLH_X1 _12285_ (.D(net276),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[13][7] ));
 DLH_X1 _12286_ (.D(net316),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[1][0] ));
 DLH_X1 _12287_ (.D(net312),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[1][1] ));
 DLH_X1 _12288_ (.D(net304),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[1][2] ));
 DLH_X1 _12289_ (.D(net298),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[1][3] ));
 DLH_X1 _12290_ (.D(net295),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[1][4] ));
 DLH_X1 _12291_ (.D(net288),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[1][5] ));
 DLH_X1 _12292_ (.D(net282),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[1][6] ));
 DLH_X1 _12293_ (.D(net276),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[1][7] ));
 DLH_X1 _12294_ (.D(net316),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[26][0] ));
 DLH_X1 _12295_ (.D(net312),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[26][1] ));
 DLH_X1 _12296_ (.D(net304),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[26][2] ));
 DLH_X1 _12297_ (.D(net298),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[26][3] ));
 DLH_X1 _12298_ (.D(net295),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[26][4] ));
 DLH_X1 _12299_ (.D(net288),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[26][5] ));
 DLH_X1 _12300_ (.D(net282),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[26][6] ));
 DLH_X1 _12301_ (.D(net276),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[26][7] ));
 DLH_X1 _12302_ (.D(net316),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[9][0] ));
 DLH_X1 _12303_ (.D(net312),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[9][1] ));
 DLH_X1 _12304_ (.D(net304),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[9][2] ));
 DLH_X1 _12305_ (.D(net298),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[9][3] ));
 DLH_X1 _12306_ (.D(net295),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[9][4] ));
 DLH_X1 _12307_ (.D(net288),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[9][5] ));
 DLH_X1 _12308_ (.D(net282),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[9][6] ));
 DLH_X1 _12309_ (.D(net276),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[9][7] ));
 DLH_X1 _12310_ (.D(net317),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[0][0] ));
 DLH_X1 _12311_ (.D(net311),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[0][1] ));
 DLH_X1 _12312_ (.D(net306),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[0][2] ));
 DLH_X1 _12313_ (.D(net300),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[0][3] ));
 DLH_X1 _12314_ (.D(net294),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[0][4] ));
 DLH_X1 _12315_ (.D(net287),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[0][5] ));
 DLH_X1 _12316_ (.D(net284),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[0][6] ));
 DLH_X1 _12317_ (.D(net277),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[0][7] ));
 DLH_X1 _12318_ (.D(net316),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[20][0] ));
 DLH_X1 _12319_ (.D(net312),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[20][1] ));
 DLH_X1 _12320_ (.D(net304),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[20][2] ));
 DLH_X1 _12321_ (.D(net298),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[20][3] ));
 DLH_X1 _12322_ (.D(net295),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[20][4] ));
 DLH_X1 _12323_ (.D(net288),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[20][5] ));
 DLH_X1 _12324_ (.D(net282),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[20][6] ));
 DLH_X1 _12325_ (.D(net276),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[20][7] ));
 DLH_X1 _12326_ (.D(net316),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[2][0] ));
 DLH_X1 _12327_ (.D(net312),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[2][1] ));
 DLH_X1 _12328_ (.D(net304),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[2][2] ));
 DLH_X1 _12329_ (.D(net298),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[2][3] ));
 DLH_X1 _12330_ (.D(net295),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[2][4] ));
 DLH_X1 _12331_ (.D(net288),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[2][5] ));
 DLH_X1 _12332_ (.D(net282),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[2][6] ));
 DLH_X1 _12333_ (.D(net276),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[2][7] ));
 DLH_X1 _12334_ (.D(net316),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[25][0] ));
 DLH_X1 _12335_ (.D(net312),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[25][1] ));
 DLH_X1 _12336_ (.D(net304),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[25][2] ));
 DLH_X1 _12337_ (.D(net298),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[25][3] ));
 DLH_X1 _12338_ (.D(net295),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[25][4] ));
 DLH_X1 _12339_ (.D(net288),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[25][5] ));
 DLH_X1 _12340_ (.D(net282),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[25][6] ));
 DLH_X1 _12341_ (.D(net276),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[25][7] ));
 DLH_X1 _12342_ (.D(net316),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[10][0] ));
 DLH_X1 _12343_ (.D(net312),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[10][1] ));
 DLH_X1 _12344_ (.D(net304),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[10][2] ));
 DLH_X1 _12345_ (.D(net298),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[10][3] ));
 DLH_X1 _12346_ (.D(net295),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[10][4] ));
 DLH_X1 _12347_ (.D(net288),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[10][5] ));
 DLH_X1 _12348_ (.D(net282),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[10][6] ));
 DLH_X1 _12349_ (.D(net276),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[10][7] ));
 DLH_X1 _12350_ (.D(net316),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[3][0] ));
 DLH_X1 _12351_ (.D(net312),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[3][1] ));
 DLH_X1 _12352_ (.D(net304),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[3][2] ));
 DLH_X1 _12353_ (.D(net298),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[3][3] ));
 DLH_X1 _12354_ (.D(net295),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[3][4] ));
 DLH_X1 _12355_ (.D(net288),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[3][5] ));
 DLH_X1 _12356_ (.D(net282),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[3][6] ));
 DLH_X1 _12357_ (.D(net276),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[3][7] ));
 DLH_X1 _12358_ (.D(net316),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[16][0] ));
 DLH_X1 _12359_ (.D(net312),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[16][1] ));
 DLH_X1 _12360_ (.D(net304),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[16][2] ));
 DLH_X1 _12361_ (.D(net298),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[16][3] ));
 DLH_X1 _12362_ (.D(net295),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[16][4] ));
 DLH_X1 _12363_ (.D(net288),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[16][5] ));
 DLH_X1 _12364_ (.D(net282),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[16][6] ));
 DLH_X1 _12365_ (.D(net276),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[16][7] ));
 DLH_X1 _12366_ (.D(net316),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[24][0] ));
 DLH_X1 _12367_ (.D(net312),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[24][1] ));
 DLH_X1 _12368_ (.D(net304),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[24][2] ));
 DLH_X1 _12369_ (.D(net298),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[24][3] ));
 DLH_X1 _12370_ (.D(net295),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[24][4] ));
 DLH_X1 _12371_ (.D(net288),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[24][5] ));
 DLH_X1 _12372_ (.D(net282),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[24][6] ));
 DLH_X1 _12373_ (.D(net276),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[24][7] ));
 DLH_X1 _12374_ (.D(net316),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[4][0] ));
 DLH_X1 _12375_ (.D(net312),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[4][1] ));
 DLH_X1 _12376_ (.D(net304),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[4][2] ));
 DLH_X1 _12377_ (.D(net298),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[4][3] ));
 DLH_X1 _12378_ (.D(net295),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[4][4] ));
 DLH_X1 _12379_ (.D(net288),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[4][5] ));
 DLH_X1 _12380_ (.D(net282),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[4][6] ));
 DLH_X1 _12381_ (.D(net276),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[4][7] ));
 DLH_X1 _12382_ (.D(net316),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[15][0] ));
 DLH_X1 _12383_ (.D(net312),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[15][1] ));
 DLH_X1 _12384_ (.D(net304),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[15][2] ));
 DLH_X1 _12385_ (.D(net298),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[15][3] ));
 DLH_X1 _12386_ (.D(net295),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[15][4] ));
 DLH_X1 _12387_ (.D(net288),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[15][5] ));
 DLH_X1 _12388_ (.D(net282),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[15][6] ));
 DLH_X1 _12389_ (.D(net276),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[15][7] ));
 DLH_X1 _12390_ (.D(net316),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[11][0] ));
 DLH_X1 _12391_ (.D(net312),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[11][1] ));
 DLH_X1 _12392_ (.D(net304),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[11][2] ));
 DLH_X1 _12393_ (.D(net298),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[11][3] ));
 DLH_X1 _12394_ (.D(net295),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[11][4] ));
 DLH_X1 _12395_ (.D(net288),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[11][5] ));
 DLH_X1 _12396_ (.D(net282),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[11][6] ));
 DLH_X1 _12397_ (.D(net276),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[11][7] ));
 DLH_X1 _12398_ (.D(net316),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[5][0] ));
 DLH_X1 _12399_ (.D(net312),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[5][1] ));
 DLH_X1 _12400_ (.D(net304),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[5][2] ));
 DLH_X1 _12401_ (.D(net298),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[5][3] ));
 DLH_X1 _12402_ (.D(net295),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[5][4] ));
 DLH_X1 _12403_ (.D(net288),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[5][5] ));
 DLH_X1 _12404_ (.D(net282),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[5][6] ));
 DLH_X1 _12405_ (.D(net276),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[5][7] ));
 DLH_X1 _12406_ (.D(net316),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[23][0] ));
 DLH_X1 _12407_ (.D(net312),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[23][1] ));
 DLH_X1 _12408_ (.D(net304),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[23][2] ));
 DLH_X1 _12409_ (.D(net298),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[23][3] ));
 DLH_X1 _12410_ (.D(net295),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[23][4] ));
 DLH_X1 _12411_ (.D(net288),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[23][5] ));
 DLH_X1 _12412_ (.D(net282),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[23][6] ));
 DLH_X1 _12413_ (.D(net276),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[23][7] ));
 DLH_X1 _12414_ (.D(net316),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[19][0] ));
 DLH_X1 _12415_ (.D(net312),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[19][1] ));
 DLH_X1 _12416_ (.D(net304),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[19][2] ));
 DLH_X1 _12417_ (.D(net298),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[19][3] ));
 DLH_X1 _12418_ (.D(net295),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[19][4] ));
 DLH_X1 _12419_ (.D(net288),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[19][5] ));
 DLH_X1 _12420_ (.D(net282),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[19][6] ));
 DLH_X1 _12421_ (.D(net276),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[19][7] ));
 DLH_X1 _12422_ (.D(net316),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[31][0] ));
 DLH_X1 _12423_ (.D(net312),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[31][1] ));
 DLH_X1 _12424_ (.D(net304),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[31][2] ));
 DLH_X1 _12425_ (.D(net298),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[31][3] ));
 DLH_X1 _12426_ (.D(net295),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[31][4] ));
 DLH_X1 _12427_ (.D(net288),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[31][5] ));
 DLH_X1 _12428_ (.D(net282),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[31][6] ));
 DLH_X1 _12429_ (.D(net276),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[31][7] ));
 DLH_X1 _12430_ (.D(net316),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[6][0] ));
 DLH_X1 _12431_ (.D(net312),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[6][1] ));
 DLH_X1 _12432_ (.D(net304),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[6][2] ));
 DLH_X1 _12433_ (.D(net298),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[6][3] ));
 DLH_X1 _12434_ (.D(net295),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[6][4] ));
 DLH_X1 _12435_ (.D(net288),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[6][5] ));
 DLH_X1 _12436_ (.D(net282),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[6][6] ));
 DLH_X1 _12437_ (.D(net276),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[6][7] ));
 DLH_X1 _12438_ (.D(net316),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[14][0] ));
 DLH_X1 _12439_ (.D(net312),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[14][1] ));
 DLH_X1 _12440_ (.D(net304),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[14][2] ));
 DLH_X1 _12441_ (.D(net298),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[14][3] ));
 DLH_X1 _12442_ (.D(net295),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[14][4] ));
 DLH_X1 _12443_ (.D(net288),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[14][5] ));
 DLH_X1 _12444_ (.D(net282),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[14][6] ));
 DLH_X1 _12445_ (.D(net276),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[14][7] ));
 DLH_X1 _12446_ (.D(net316),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[30][0] ));
 DLH_X1 _12447_ (.D(net312),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[30][1] ));
 DLH_X1 _12448_ (.D(net304),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[30][2] ));
 DLH_X1 _12449_ (.D(net298),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[30][3] ));
 DLH_X1 _12450_ (.D(net295),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[30][4] ));
 DLH_X1 _12451_ (.D(net288),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[30][5] ));
 DLH_X1 _12452_ (.D(net282),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[30][6] ));
 DLH_X1 _12453_ (.D(net276),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[30][7] ));
 DLH_X1 _12454_ (.D(net316),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[22][0] ));
 DLH_X1 _12455_ (.D(net312),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[22][1] ));
 DLH_X1 _12456_ (.D(net304),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[22][2] ));
 DLH_X1 _12457_ (.D(net298),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[22][3] ));
 DLH_X1 _12458_ (.D(net295),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[22][4] ));
 DLH_X1 _12459_ (.D(net288),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[22][5] ));
 DLH_X1 _12460_ (.D(net282),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[22][6] ));
 DLH_X1 _12461_ (.D(net276),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[22][7] ));
 DLH_X1 _12462_ (.D(net316),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[7][0] ));
 DLH_X1 _12463_ (.D(net312),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[7][1] ));
 DLH_X1 _12464_ (.D(net304),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[7][2] ));
 DLH_X1 _12465_ (.D(net298),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[7][3] ));
 DLH_X1 _12466_ (.D(net295),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[7][4] ));
 DLH_X1 _12467_ (.D(net288),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[7][5] ));
 DLH_X1 _12468_ (.D(net282),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[7][6] ));
 DLH_X1 _12469_ (.D(net276),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[7][7] ));
 DLH_X1 _12470_ (.D(net316),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[29][0] ));
 DLH_X1 _12471_ (.D(net312),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[29][1] ));
 DLH_X1 _12472_ (.D(net304),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[29][2] ));
 DLH_X1 _12473_ (.D(net298),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[29][3] ));
 DLH_X1 _12474_ (.D(net295),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[29][4] ));
 DLH_X1 _12475_ (.D(net288),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[29][5] ));
 DLH_X1 _12476_ (.D(net282),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[29][6] ));
 DLH_X1 _12477_ (.D(net276),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[29][7] ));
 DLH_X1 _12478_ (.D(net316),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[12][0] ));
 DLH_X1 _12479_ (.D(net312),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[12][1] ));
 DLH_X1 _12480_ (.D(net304),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[12][2] ));
 DLH_X1 _12481_ (.D(net298),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[12][3] ));
 DLH_X1 _12482_ (.D(net295),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[12][4] ));
 DLH_X1 _12483_ (.D(net288),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[12][5] ));
 DLH_X1 _12484_ (.D(net282),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[12][6] ));
 DLH_X1 _12485_ (.D(net276),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[12][7] ));
 DLH_X1 _12486_ (.D(net316),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[17][0] ));
 DLH_X1 _12487_ (.D(net312),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[17][1] ));
 DLH_X1 _12488_ (.D(net304),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[17][2] ));
 DLH_X1 _12489_ (.D(net298),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[17][3] ));
 DLH_X1 _12490_ (.D(net295),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[17][4] ));
 DLH_X1 _12491_ (.D(net288),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[17][5] ));
 DLH_X1 _12492_ (.D(net282),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[17][6] ));
 DLH_X1 _12493_ (.D(net276),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[17][7] ));
 DLH_X1 _12494_ (.D(net316),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[28][0] ));
 DLH_X1 _12495_ (.D(net312),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[28][1] ));
 DLH_X1 _12496_ (.D(net304),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[28][2] ));
 DLH_X1 _12497_ (.D(net298),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[28][3] ));
 DLH_X1 _12498_ (.D(net295),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[28][4] ));
 DLH_X1 _12499_ (.D(net288),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[28][5] ));
 DLH_X1 _12500_ (.D(net282),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[28][6] ));
 DLH_X1 _12501_ (.D(net276),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[28][7] ));
 DLH_X1 _12502_ (.D(net316),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[8][0] ));
 DLH_X1 _12503_ (.D(net312),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[8][1] ));
 DLH_X1 _12504_ (.D(net304),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[8][2] ));
 DLH_X1 _12505_ (.D(net298),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[8][3] ));
 DLH_X1 _12506_ (.D(net295),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[8][4] ));
 DLH_X1 _12507_ (.D(net288),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[8][5] ));
 DLH_X1 _12508_ (.D(net282),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[8][6] ));
 DLH_X1 _12509_ (.D(net276),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[8][7] ));
 DLH_X1 _12510_ (.D(net316),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[21][0] ));
 DLH_X1 _12511_ (.D(net312),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[21][1] ));
 DLH_X1 _12512_ (.D(net304),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[21][2] ));
 DLH_X1 _12513_ (.D(net298),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[21][3] ));
 DLH_X1 _12514_ (.D(net295),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[21][4] ));
 DLH_X1 _12515_ (.D(net288),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[21][5] ));
 DLH_X1 _12516_ (.D(net282),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[21][6] ));
 DLH_X1 _12517_ (.D(net276),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[21][7] ));
 DLH_X1 _12518_ (.D(net316),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[27][0] ));
 DLH_X1 _12519_ (.D(net312),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[27][1] ));
 DLH_X1 _12520_ (.D(net304),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[27][2] ));
 DLH_X1 _12521_ (.D(net298),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[27][3] ));
 DLH_X1 _12522_ (.D(net295),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[27][4] ));
 DLH_X1 _12523_ (.D(net288),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[27][5] ));
 DLH_X1 _12524_ (.D(net282),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[27][6] ));
 DLH_X1 _12525_ (.D(net276),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[27][7] ));
 DLH_X1 _12526_ (.D(net316),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[18][0] ));
 DLH_X1 _12527_ (.D(net312),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[18][1] ));
 DLH_X1 _12528_ (.D(net304),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[18][2] ));
 DLH_X1 _12529_ (.D(net298),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[18][3] ));
 DLH_X1 _12530_ (.D(net295),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[18][4] ));
 DLH_X1 _12531_ (.D(net288),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[18][5] ));
 DLH_X1 _12532_ (.D(net282),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[18][6] ));
 DLH_X1 _12533_ (.D(net276),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.mem[18][7] ));
 DLL_X1 _12534_ (.D(\lut.gen_sub_units_scm.__6.sub_unit_i.cg_we_global.en_i ),
    .GN(clknet_level_5_1_114__00532_),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.cg_we_global.clk_en ));
 DLL_X1 _12535_ (.D(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__0.cg_i.en_i ),
    .GN(clknet_level_2_1_498__00561_),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_en ));
 DLL_X1 _12536_ (.D(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__1.cg_i.en_i ),
    .GN(clknet_level_2_1_292__00561_),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_en ));
 DLL_X1 _12537_ (.D(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__2.cg_i.en_i ),
    .GN(clknet_level_2_1_498__00561_),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_en ));
 DLL_X1 _12538_ (.D(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__3.cg_i.en_i ),
    .GN(clknet_level_2_1_5101__00561_),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_en ));
 DLL_X1 _12539_ (.D(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__4.cg_i.en_i ),
    .GN(clknet_level_2_1_395__00561_),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_en ));
 DLL_X1 _12540_ (.D(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__5.cg_i.en_i ),
    .GN(clknet_level_2_1_292__00561_),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_en ));
 DLL_X1 _12541_ (.D(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__6.cg_i.en_i ),
    .GN(clknet_level_2_1_8110__00561_),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_en ));
 DLL_X1 _12542_ (.D(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__7.cg_i.en_i ),
    .GN(clknet_level_2_1_498__00561_),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_en ));
 DLL_X1 _12543_ (.D(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__8.cg_i.en_i ),
    .GN(clknet_level_2_1_395__00561_),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_en ));
 DLL_X1 _12544_ (.D(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__9.cg_i.en_i ),
    .GN(clknet_level_2_1_395__00561_),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_en ));
 DLL_X1 _12545_ (.D(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__10.cg_i.en_i ),
    .GN(clknet_level_2_1_189__00561_),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_en ));
 DLL_X1 _12546_ (.D(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__11.cg_i.en_i ),
    .GN(clknet_level_2_1_8110__00561_),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_en ));
 DLL_X1 _12547_ (.D(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__12.cg_i.en_i ),
    .GN(clknet_level_2_1_498__00561_),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_en ));
 DLL_X1 _12548_ (.D(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__13.cg_i.en_i ),
    .GN(clknet_level_2_1_292__00561_),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_en ));
 DLL_X1 _12549_ (.D(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__14.cg_i.en_i ),
    .GN(clknet_level_2_1_8110__00561_),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_en ));
 DLL_X1 _12550_ (.D(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__15.cg_i.en_i ),
    .GN(clknet_level_2_1_5101__00561_),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_en ));
 DLL_X1 _12551_ (.D(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__16.cg_i.en_i ),
    .GN(clknet_level_2_1_6104__00561_),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_en ));
 DLL_X1 _12552_ (.D(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__17.cg_i.en_i ),
    .GN(clknet_level_2_1_5101__00561_),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_en ));
 DLL_X1 _12553_ (.D(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__18.cg_i.en_i ),
    .GN(clknet_level_2_1_189__00561_),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_en ));
 DLL_X1 _12554_ (.D(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__19.cg_i.en_i ),
    .GN(clknet_level_2_1_189__00561_),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_en ));
 DLL_X1 _12555_ (.D(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__20.cg_i.en_i ),
    .GN(clknet_level_2_1_5101__00561_),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_en ));
 DLL_X1 _12556_ (.D(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__21.cg_i.en_i ),
    .GN(clknet_level_2_1_6104__00561_),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_en ));
 DLL_X1 _12557_ (.D(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__22.cg_i.en_i ),
    .GN(clknet_level_2_1_395__00561_),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_en ));
 DLL_X1 _12558_ (.D(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__23.cg_i.en_i ),
    .GN(clknet_level_2_1_5101__00561_),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_en ));
 DLL_X1 _12559_ (.D(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__24.cg_i.en_i ),
    .GN(clknet_level_2_1_7107__00561_),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_en ));
 DLL_X1 _12560_ (.D(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__25.cg_i.en_i ),
    .GN(clknet_level_2_1_189__00561_),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_en ));
 DLL_X1 _12561_ (.D(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__26.cg_i.en_i ),
    .GN(clknet_level_2_1_189__00561_),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_en ));
 DLL_X1 _12562_ (.D(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__27.cg_i.en_i ),
    .GN(clknet_level_2_1_7107__00561_),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_en ));
 DLL_X1 _12563_ (.D(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__28.cg_i.en_i ),
    .GN(clknet_level_2_1_395__00561_),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_en ));
 DLL_X1 _12564_ (.D(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__29.cg_i.en_i ),
    .GN(clknet_level_2_1_292__00561_),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_en ));
 DLL_X1 _12565_ (.D(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__30.cg_i.en_i ),
    .GN(clknet_level_2_1_395__00561_),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_en ));
 DLL_X1 _12566_ (.D(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__31.cg_i.en_i ),
    .GN(clknet_level_2_1_189__00561_),
    .Q(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_en ));
 DLH_X1 _12567_ (.D(net321),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[13][0] ));
 DLH_X1 _12568_ (.D(net310),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[13][1] ));
 DLH_X1 _12569_ (.D(net308),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[13][2] ));
 DLH_X1 _12570_ (.D(net302),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[13][3] ));
 DLH_X1 _12571_ (.D(net293),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[13][4] ));
 DLH_X1 _12572_ (.D(net291),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[13][5] ));
 DLH_X1 _12573_ (.D(net283),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[13][6] ));
 DLH_X1 _12574_ (.D(net280),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[13][7] ));
 DLH_X1 _12575_ (.D(net321),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[1][0] ));
 DLH_X1 _12576_ (.D(net310),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[1][1] ));
 DLH_X1 _12577_ (.D(net308),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[1][2] ));
 DLH_X1 _12578_ (.D(net302),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[1][3] ));
 DLH_X1 _12579_ (.D(net297),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[1][4] ));
 DLH_X1 _12580_ (.D(net291),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[1][5] ));
 DLH_X1 _12581_ (.D(net283),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[1][6] ));
 DLH_X1 _12582_ (.D(net280),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[1][7] ));
 DLH_X1 _12583_ (.D(net321),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[26][0] ));
 DLH_X1 _12584_ (.D(net310),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[26][1] ));
 DLH_X1 _12585_ (.D(net308),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[26][2] ));
 DLH_X1 _12586_ (.D(net300),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[26][3] ));
 DLH_X1 _12587_ (.D(net297),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[26][4] ));
 DLH_X1 _12588_ (.D(net291),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[26][5] ));
 DLH_X1 _12589_ (.D(net283),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[26][6] ));
 DLH_X1 _12590_ (.D(net280),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[26][7] ));
 DLH_X1 _12591_ (.D(net321),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[9][0] ));
 DLH_X1 _12592_ (.D(net310),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[9][1] ));
 DLH_X1 _12593_ (.D(net308),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[9][2] ));
 DLH_X1 _12594_ (.D(net300),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[9][3] ));
 DLH_X1 _12595_ (.D(net293),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[9][4] ));
 DLH_X1 _12596_ (.D(net291),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[9][5] ));
 DLH_X1 _12597_ (.D(net283),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[9][6] ));
 DLH_X1 _12598_ (.D(net280),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[9][7] ));
 DLH_X1 _12599_ (.D(net319),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[0][0] ));
 DLH_X1 _12600_ (.D(net311),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[0][1] ));
 DLH_X1 _12601_ (.D(net305),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[0][2] ));
 DLH_X1 _12602_ (.D(net300),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[0][3] ));
 DLH_X1 _12603_ (.D(net294),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[0][4] ));
 DLH_X1 _12604_ (.D(net287),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[0][5] ));
 DLH_X1 _12605_ (.D(net285),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[0][6] ));
 DLH_X1 _12606_ (.D(net277),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[0][7] ));
 DLH_X1 _12607_ (.D(net321),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[20][0] ));
 DLH_X1 _12608_ (.D(net310),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[20][1] ));
 DLH_X1 _12609_ (.D(net308),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[20][2] ));
 DLH_X1 _12610_ (.D(net302),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[20][3] ));
 DLH_X1 _12611_ (.D(net297),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[20][4] ));
 DLH_X1 _12612_ (.D(net291),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[20][5] ));
 DLH_X1 _12613_ (.D(net283),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[20][6] ));
 DLH_X1 _12614_ (.D(net280),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[20][7] ));
 DLH_X1 _12615_ (.D(net321),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[2][0] ));
 DLH_X1 _12616_ (.D(net310),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[2][1] ));
 DLH_X1 _12617_ (.D(net308),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[2][2] ));
 DLH_X1 _12618_ (.D(net302),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[2][3] ));
 DLH_X1 _12619_ (.D(net293),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[2][4] ));
 DLH_X1 _12620_ (.D(net291),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[2][5] ));
 DLH_X1 _12621_ (.D(net283),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[2][6] ));
 DLH_X1 _12622_ (.D(net280),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[2][7] ));
 DLH_X1 _12623_ (.D(net321),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[25][0] ));
 DLH_X1 _12624_ (.D(net310),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[25][1] ));
 DLH_X1 _12625_ (.D(net308),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[25][2] ));
 DLH_X1 _12626_ (.D(net302),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[25][3] ));
 DLH_X1 _12627_ (.D(net293),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[25][4] ));
 DLH_X1 _12628_ (.D(net291),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[25][5] ));
 DLH_X1 _12629_ (.D(net283),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[25][6] ));
 DLH_X1 _12630_ (.D(net280),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[25][7] ));
 DLH_X1 _12631_ (.D(net321),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[10][0] ));
 DLH_X1 _12632_ (.D(net310),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[10][1] ));
 DLH_X1 _12633_ (.D(net308),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[10][2] ));
 DLH_X1 _12634_ (.D(net300),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[10][3] ));
 DLH_X1 _12635_ (.D(net297),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[10][4] ));
 DLH_X1 _12636_ (.D(net291),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[10][5] ));
 DLH_X1 _12637_ (.D(net283),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[10][6] ));
 DLH_X1 _12638_ (.D(net280),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[10][7] ));
 DLH_X1 _12639_ (.D(net321),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[3][0] ));
 DLH_X1 _12640_ (.D(net310),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[3][1] ));
 DLH_X1 _12641_ (.D(net308),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[3][2] ));
 DLH_X1 _12642_ (.D(net300),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[3][3] ));
 DLH_X1 _12643_ (.D(net297),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[3][4] ));
 DLH_X1 _12644_ (.D(net291),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[3][5] ));
 DLH_X1 _12645_ (.D(net283),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[3][6] ));
 DLH_X1 _12646_ (.D(net280),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[3][7] ));
 DLH_X1 _12647_ (.D(net321),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[16][0] ));
 DLH_X1 _12648_ (.D(net310),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[16][1] ));
 DLH_X1 _12649_ (.D(net308),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[16][2] ));
 DLH_X1 _12650_ (.D(net302),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[16][3] ));
 DLH_X1 _12651_ (.D(net297),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[16][4] ));
 DLH_X1 _12652_ (.D(net291),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[16][5] ));
 DLH_X1 _12653_ (.D(net283),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[16][6] ));
 DLH_X1 _12654_ (.D(net280),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[16][7] ));
 DLH_X1 _12655_ (.D(net321),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[24][0] ));
 DLH_X1 _12656_ (.D(net310),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[24][1] ));
 DLH_X1 _12657_ (.D(net308),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[24][2] ));
 DLH_X1 _12658_ (.D(net300),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[24][3] ));
 DLH_X1 _12659_ (.D(net297),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[24][4] ));
 DLH_X1 _12660_ (.D(net291),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[24][5] ));
 DLH_X1 _12661_ (.D(net283),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[24][6] ));
 DLH_X1 _12662_ (.D(net280),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[24][7] ));
 DLH_X1 _12663_ (.D(net321),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[4][0] ));
 DLH_X1 _12664_ (.D(net310),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[4][1] ));
 DLH_X1 _12665_ (.D(net308),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[4][2] ));
 DLH_X1 _12666_ (.D(net300),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[4][3] ));
 DLH_X1 _12667_ (.D(net297),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[4][4] ));
 DLH_X1 _12668_ (.D(net291),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[4][5] ));
 DLH_X1 _12669_ (.D(net283),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[4][6] ));
 DLH_X1 _12670_ (.D(net280),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[4][7] ));
 DLH_X1 _12671_ (.D(net321),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[15][0] ));
 DLH_X1 _12672_ (.D(net310),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[15][1] ));
 DLH_X1 _12673_ (.D(net308),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[15][2] ));
 DLH_X1 _12674_ (.D(net302),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[15][3] ));
 DLH_X1 _12675_ (.D(net293),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[15][4] ));
 DLH_X1 _12676_ (.D(net291),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[15][5] ));
 DLH_X1 _12677_ (.D(net283),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[15][6] ));
 DLH_X1 _12678_ (.D(net280),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[15][7] ));
 DLH_X1 _12679_ (.D(net321),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[11][0] ));
 DLH_X1 _12680_ (.D(net310),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[11][1] ));
 DLH_X1 _12681_ (.D(net308),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[11][2] ));
 DLH_X1 _12682_ (.D(net302),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[11][3] ));
 DLH_X1 _12683_ (.D(net293),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[11][4] ));
 DLH_X1 _12684_ (.D(net291),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[11][5] ));
 DLH_X1 _12685_ (.D(net283),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[11][6] ));
 DLH_X1 _12686_ (.D(net280),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[11][7] ));
 DLH_X1 _12687_ (.D(net321),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[5][0] ));
 DLH_X1 _12688_ (.D(net310),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[5][1] ));
 DLH_X1 _12689_ (.D(net308),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[5][2] ));
 DLH_X1 _12690_ (.D(net302),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[5][3] ));
 DLH_X1 _12691_ (.D(net297),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[5][4] ));
 DLH_X1 _12692_ (.D(net291),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[5][5] ));
 DLH_X1 _12693_ (.D(net283),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[5][6] ));
 DLH_X1 _12694_ (.D(net280),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[5][7] ));
 DLH_X1 _12695_ (.D(net321),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[23][0] ));
 DLH_X1 _12696_ (.D(net310),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[23][1] ));
 DLH_X1 _12697_ (.D(net308),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[23][2] ));
 DLH_X1 _12698_ (.D(net302),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[23][3] ));
 DLH_X1 _12699_ (.D(net297),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[23][4] ));
 DLH_X1 _12700_ (.D(net291),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[23][5] ));
 DLH_X1 _12701_ (.D(net283),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[23][6] ));
 DLH_X1 _12702_ (.D(net280),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[23][7] ));
 DLH_X1 _12703_ (.D(net321),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[19][0] ));
 DLH_X1 _12704_ (.D(net310),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[19][1] ));
 DLH_X1 _12705_ (.D(net308),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[19][2] ));
 DLH_X1 _12706_ (.D(net302),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[19][3] ));
 DLH_X1 _12707_ (.D(net297),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[19][4] ));
 DLH_X1 _12708_ (.D(net291),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[19][5] ));
 DLH_X1 _12709_ (.D(net283),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[19][6] ));
 DLH_X1 _12710_ (.D(net280),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[19][7] ));
 DLH_X1 _12711_ (.D(net321),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[31][0] ));
 DLH_X1 _12712_ (.D(net310),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[31][1] ));
 DLH_X1 _12713_ (.D(net308),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[31][2] ));
 DLH_X1 _12714_ (.D(net300),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[31][3] ));
 DLH_X1 _12715_ (.D(net297),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[31][4] ));
 DLH_X1 _12716_ (.D(net291),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[31][5] ));
 DLH_X1 _12717_ (.D(net283),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[31][6] ));
 DLH_X1 _12718_ (.D(net280),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[31][7] ));
 DLH_X1 _12719_ (.D(net321),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[6][0] ));
 DLH_X1 _12720_ (.D(net310),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[6][1] ));
 DLH_X1 _12721_ (.D(net308),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[6][2] ));
 DLH_X1 _12722_ (.D(net302),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[6][3] ));
 DLH_X1 _12723_ (.D(net297),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[6][4] ));
 DLH_X1 _12724_ (.D(net291),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[6][5] ));
 DLH_X1 _12725_ (.D(net283),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[6][6] ));
 DLH_X1 _12726_ (.D(net280),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[6][7] ));
 DLH_X1 _12727_ (.D(net321),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[14][0] ));
 DLH_X1 _12728_ (.D(net310),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[14][1] ));
 DLH_X1 _12729_ (.D(net308),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[14][2] ));
 DLH_X1 _12730_ (.D(net300),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[14][3] ));
 DLH_X1 _12731_ (.D(net293),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[14][4] ));
 DLH_X1 _12732_ (.D(net291),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[14][5] ));
 DLH_X1 _12733_ (.D(net283),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[14][6] ));
 DLH_X1 _12734_ (.D(net280),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[14][7] ));
 DLH_X1 _12735_ (.D(net321),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[30][0] ));
 DLH_X1 _12736_ (.D(net310),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[30][1] ));
 DLH_X1 _12737_ (.D(net308),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[30][2] ));
 DLH_X1 _12738_ (.D(net302),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[30][3] ));
 DLH_X1 _12739_ (.D(net293),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[30][4] ));
 DLH_X1 _12740_ (.D(net291),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[30][5] ));
 DLH_X1 _12741_ (.D(net283),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[30][6] ));
 DLH_X1 _12742_ (.D(net280),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[30][7] ));
 DLH_X1 _12743_ (.D(net321),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[22][0] ));
 DLH_X1 _12744_ (.D(net310),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[22][1] ));
 DLH_X1 _12745_ (.D(net308),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[22][2] ));
 DLH_X1 _12746_ (.D(net300),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[22][3] ));
 DLH_X1 _12747_ (.D(net293),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[22][4] ));
 DLH_X1 _12748_ (.D(net291),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[22][5] ));
 DLH_X1 _12749_ (.D(net283),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[22][6] ));
 DLH_X1 _12750_ (.D(net280),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[22][7] ));
 DLH_X1 _12751_ (.D(net321),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[7][0] ));
 DLH_X1 _12752_ (.D(net310),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[7][1] ));
 DLH_X1 _12753_ (.D(net308),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[7][2] ));
 DLH_X1 _12754_ (.D(net302),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[7][3] ));
 DLH_X1 _12755_ (.D(net297),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[7][4] ));
 DLH_X1 _12756_ (.D(net291),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[7][5] ));
 DLH_X1 _12757_ (.D(net283),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[7][6] ));
 DLH_X1 _12758_ (.D(net280),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[7][7] ));
 DLH_X1 _12759_ (.D(net321),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[29][0] ));
 DLH_X1 _12760_ (.D(net310),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[29][1] ));
 DLH_X1 _12761_ (.D(net308),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[29][2] ));
 DLH_X1 _12762_ (.D(net300),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[29][3] ));
 DLH_X1 _12763_ (.D(net297),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[29][4] ));
 DLH_X1 _12764_ (.D(net291),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[29][5] ));
 DLH_X1 _12765_ (.D(net283),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[29][6] ));
 DLH_X1 _12766_ (.D(net280),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[29][7] ));
 DLH_X1 _12767_ (.D(net321),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[12][0] ));
 DLH_X1 _12768_ (.D(net310),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[12][1] ));
 DLH_X1 _12769_ (.D(net308),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[12][2] ));
 DLH_X1 _12770_ (.D(net300),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[12][3] ));
 DLH_X1 _12771_ (.D(net293),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[12][4] ));
 DLH_X1 _12772_ (.D(net291),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[12][5] ));
 DLH_X1 _12773_ (.D(net283),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[12][6] ));
 DLH_X1 _12774_ (.D(net280),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[12][7] ));
 DLH_X1 _12775_ (.D(net321),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[17][0] ));
 DLH_X1 _12776_ (.D(net310),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[17][1] ));
 DLH_X1 _12777_ (.D(net308),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[17][2] ));
 DLH_X1 _12778_ (.D(net300),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[17][3] ));
 DLH_X1 _12779_ (.D(net293),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[17][4] ));
 DLH_X1 _12780_ (.D(net291),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[17][5] ));
 DLH_X1 _12781_ (.D(net283),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[17][6] ));
 DLH_X1 _12782_ (.D(net280),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[17][7] ));
 DLH_X1 _12783_ (.D(net321),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[28][0] ));
 DLH_X1 _12784_ (.D(net310),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[28][1] ));
 DLH_X1 _12785_ (.D(net308),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[28][2] ));
 DLH_X1 _12786_ (.D(net300),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[28][3] ));
 DLH_X1 _12787_ (.D(net297),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[28][4] ));
 DLH_X1 _12788_ (.D(net291),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[28][5] ));
 DLH_X1 _12789_ (.D(net283),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[28][6] ));
 DLH_X1 _12790_ (.D(net280),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[28][7] ));
 DLH_X1 _12791_ (.D(net321),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[8][0] ));
 DLH_X1 _12792_ (.D(net310),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[8][1] ));
 DLH_X1 _12793_ (.D(net308),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[8][2] ));
 DLH_X1 _12794_ (.D(net302),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[8][3] ));
 DLH_X1 _12795_ (.D(net297),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[8][4] ));
 DLH_X1 _12796_ (.D(net291),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[8][5] ));
 DLH_X1 _12797_ (.D(net283),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[8][6] ));
 DLH_X1 _12798_ (.D(net280),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[8][7] ));
 DLH_X1 _12799_ (.D(net321),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[21][0] ));
 DLH_X1 _12800_ (.D(net310),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[21][1] ));
 DLH_X1 _12801_ (.D(net308),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[21][2] ));
 DLH_X1 _12802_ (.D(net302),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[21][3] ));
 DLH_X1 _12803_ (.D(net297),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[21][4] ));
 DLH_X1 _12804_ (.D(net291),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[21][5] ));
 DLH_X1 _12805_ (.D(net283),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[21][6] ));
 DLH_X1 _12806_ (.D(net280),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[21][7] ));
 DLH_X1 _12807_ (.D(net321),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[27][0] ));
 DLH_X1 _12808_ (.D(net310),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[27][1] ));
 DLH_X1 _12809_ (.D(net308),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[27][2] ));
 DLH_X1 _12810_ (.D(net300),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[27][3] ));
 DLH_X1 _12811_ (.D(net297),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[27][4] ));
 DLH_X1 _12812_ (.D(net291),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[27][5] ));
 DLH_X1 _12813_ (.D(net283),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[27][6] ));
 DLH_X1 _12814_ (.D(net280),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[27][7] ));
 DLH_X1 _12815_ (.D(net321),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[18][0] ));
 DLH_X1 _12816_ (.D(net310),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[18][1] ));
 DLH_X1 _12817_ (.D(net308),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[18][2] ));
 DLH_X1 _12818_ (.D(net300),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[18][3] ));
 DLH_X1 _12819_ (.D(net297),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[18][4] ));
 DLH_X1 _12820_ (.D(net291),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[18][5] ));
 DLH_X1 _12821_ (.D(net283),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[18][6] ));
 DLH_X1 _12822_ (.D(net280),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.mem[18][7] ));
 DLL_X1 _12823_ (.D(\lut.gen_sub_units_scm.__5.sub_unit_i.cg_we_global.en_i ),
    .GN(clknet_level_5_1_3218__00532_),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.cg_we_global.clk_en ));
 DLL_X1 _12824_ (.D(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__0.cg_i.en_i ),
    .GN(clknet_level_2_1_2248__00564_),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_en ));
 DLL_X1 _12825_ (.D(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__1.cg_i.en_i ),
    .GN(clknet_level_2_1_6260__00564_),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_en ));
 DLL_X1 _12826_ (.D(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__2.cg_i.en_i ),
    .GN(clknet_level_2_1_3251__00564_),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_en ));
 DLL_X1 _12827_ (.D(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__3.cg_i.en_i ),
    .GN(clknet_level_2_1_2248__00564_),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_en ));
 DLL_X1 _12828_ (.D(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__4.cg_i.en_i ),
    .GN(clknet_level_2_1_1245__00564_),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_en ));
 DLL_X1 _12829_ (.D(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__5.cg_i.en_i ),
    .GN(clknet_level_2_1_3251__00564_),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_en ));
 DLL_X1 _12830_ (.D(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__6.cg_i.en_i ),
    .GN(clknet_level_2_1_5257__00564_),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_en ));
 DLL_X1 _12831_ (.D(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__7.cg_i.en_i ),
    .GN(clknet_level_2_1_8266__00564_),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_en ));
 DLL_X1 _12832_ (.D(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__8.cg_i.en_i ),
    .GN(clknet_level_2_1_2248__00564_),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_en ));
 DLL_X1 _12833_ (.D(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__9.cg_i.en_i ),
    .GN(clknet_level_2_1_4254__00564_),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_en ));
 DLL_X1 _12834_ (.D(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__10.cg_i.en_i ),
    .GN(clknet_level_2_1_2248__00564_),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_en ));
 DLL_X1 _12835_ (.D(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__11.cg_i.en_i ),
    .GN(clknet_level_2_1_4254__00564_),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_en ));
 DLL_X1 _12836_ (.D(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__12.cg_i.en_i ),
    .GN(clknet_level_2_1_3251__00564_),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_en ));
 DLL_X1 _12837_ (.D(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__13.cg_i.en_i ),
    .GN(clknet_level_2_1_1245__00564_),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_en ));
 DLL_X1 _12838_ (.D(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__14.cg_i.en_i ),
    .GN(clknet_level_2_1_4254__00564_),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_en ));
 DLL_X1 _12839_ (.D(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__15.cg_i.en_i ),
    .GN(clknet_level_2_1_4254__00564_),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_en ));
 DLL_X1 _12840_ (.D(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__16.cg_i.en_i ),
    .GN(clknet_level_2_1_5257__00564_),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_en ));
 DLL_X1 _12841_ (.D(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__17.cg_i.en_i ),
    .GN(clknet_level_2_1_4254__00564_),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_en ));
 DLL_X1 _12842_ (.D(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__18.cg_i.en_i ),
    .GN(clknet_level_2_1_1245__00564_),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_en ));
 DLL_X1 _12843_ (.D(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__19.cg_i.en_i ),
    .GN(clknet_level_2_1_8266__00564_),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_en ));
 DLL_X1 _12844_ (.D(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__20.cg_i.en_i ),
    .GN(clknet_level_2_1_7263__00564_),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_en ));
 DLL_X1 _12845_ (.D(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__21.cg_i.en_i ),
    .GN(clknet_level_2_1_3251__00564_),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_en ));
 DLL_X1 _12846_ (.D(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__22.cg_i.en_i ),
    .GN(clknet_level_2_1_1245__00564_),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_en ));
 DLL_X1 _12847_ (.D(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__23.cg_i.en_i ),
    .GN(clknet_level_2_1_8266__00564_),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_en ));
 DLL_X1 _12848_ (.D(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__24.cg_i.en_i ),
    .GN(clknet_level_2_1_6260__00564_),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_en ));
 DLL_X1 _12849_ (.D(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__25.cg_i.en_i ),
    .GN(clknet_level_2_1_7263__00564_),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_en ));
 DLL_X1 _12850_ (.D(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__26.cg_i.en_i ),
    .GN(clknet_level_2_1_8266__00564_),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_en ));
 DLL_X1 _12851_ (.D(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__27.cg_i.en_i ),
    .GN(clknet_level_2_1_1245__00564_),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_en ));
 DLL_X1 _12852_ (.D(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__28.cg_i.en_i ),
    .GN(clknet_level_2_1_1245__00564_),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_en ));
 DLL_X1 _12853_ (.D(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__29.cg_i.en_i ),
    .GN(clknet_level_2_1_8266__00564_),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_en ));
 DLL_X1 _12854_ (.D(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__30.cg_i.en_i ),
    .GN(clknet_level_2_1_4254__00564_),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_en ));
 DLL_X1 _12855_ (.D(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__31.cg_i.en_i ),
    .GN(clknet_level_2_1_6260__00564_),
    .Q(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_en ));
 DLH_X1 _12856_ (.D(net319),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[13][0] ));
 DLH_X1 _12857_ (.D(net314),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[13][1] ));
 DLH_X1 _12858_ (.D(net309),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[13][2] ));
 DLH_X1 _12859_ (.D(net301),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[13][3] ));
 DLH_X1 _12860_ (.D(net296),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[13][4] ));
 DLH_X1 _12861_ (.D(net290),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[13][5] ));
 DLH_X1 _12862_ (.D(net286),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[13][6] ));
 DLH_X1 _12863_ (.D(net278),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[13][7] ));
 DLH_X1 _12864_ (.D(net318),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[1][0] ));
 DLH_X1 _12865_ (.D(net314),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[1][1] ));
 DLH_X1 _12866_ (.D(net307),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[1][2] ));
 DLH_X1 _12867_ (.D(net301),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[1][3] ));
 DLH_X1 _12868_ (.D(net296),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[1][4] ));
 DLH_X1 _12869_ (.D(net290),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[1][5] ));
 DLH_X1 _12870_ (.D(net281),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[1][6] ));
 DLH_X1 _12871_ (.D(net279),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[1][7] ));
 DLH_X1 _12872_ (.D(net318),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[26][0] ));
 DLH_X1 _12873_ (.D(net314),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[26][1] ));
 DLH_X1 _12874_ (.D(net307),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[26][2] ));
 DLH_X1 _12875_ (.D(net301),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[26][3] ));
 DLH_X1 _12876_ (.D(net296),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[26][4] ));
 DLH_X1 _12877_ (.D(net289),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[26][5] ));
 DLH_X1 _12878_ (.D(net281),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[26][6] ));
 DLH_X1 _12879_ (.D(net278),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[26][7] ));
 DLH_X1 _12880_ (.D(net318),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[9][0] ));
 DLH_X1 _12881_ (.D(net314),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[9][1] ));
 DLH_X1 _12882_ (.D(net309),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[9][2] ));
 DLH_X1 _12883_ (.D(net301),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[9][3] ));
 DLH_X1 _12884_ (.D(net296),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[9][4] ));
 DLH_X1 _12885_ (.D(net290),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[9][5] ));
 DLH_X1 _12886_ (.D(net286),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[9][6] ));
 DLH_X1 _12887_ (.D(net278),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[9][7] ));
 DLH_X1 _12888_ (.D(net319),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[0][0] ));
 DLH_X1 _12889_ (.D(net313),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[0][1] ));
 DLH_X1 _12890_ (.D(net306),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[0][2] ));
 DLH_X1 _12891_ (.D(net303),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[0][3] ));
 DLH_X1 _12892_ (.D(net295),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[0][4] ));
 DLH_X1 _12893_ (.D(net292),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[0][5] ));
 DLH_X1 _12894_ (.D(net285),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[0][6] ));
 DLH_X1 _12895_ (.D(net279),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[0][7] ));
 DLH_X1 _12896_ (.D(net319),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[20][0] ));
 DLH_X1 _12897_ (.D(net314),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[20][1] ));
 DLH_X1 _12898_ (.D(net309),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[20][2] ));
 DLH_X1 _12899_ (.D(net301),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[20][3] ));
 DLH_X1 _12900_ (.D(net296),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[20][4] ));
 DLH_X1 _12901_ (.D(net290),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[20][5] ));
 DLH_X1 _12902_ (.D(net286),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[20][6] ));
 DLH_X1 _12903_ (.D(net278),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[20][7] ));
 DLH_X1 _12904_ (.D(net318),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[2][0] ));
 DLH_X1 _12905_ (.D(net314),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[2][1] ));
 DLH_X1 _12906_ (.D(net307),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[2][2] ));
 DLH_X1 _12907_ (.D(net301),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[2][3] ));
 DLH_X1 _12908_ (.D(net296),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[2][4] ));
 DLH_X1 _12909_ (.D(net290),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[2][5] ));
 DLH_X1 _12910_ (.D(net281),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[2][6] ));
 DLH_X1 _12911_ (.D(net278),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[2][7] ));
 DLH_X1 _12912_ (.D(net319),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[25][0] ));
 DLH_X1 _12913_ (.D(net314),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[25][1] ));
 DLH_X1 _12914_ (.D(net309),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[25][2] ));
 DLH_X1 _12915_ (.D(net301),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[25][3] ));
 DLH_X1 _12916_ (.D(net296),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[25][4] ));
 DLH_X1 _12917_ (.D(net290),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[25][5] ));
 DLH_X1 _12918_ (.D(net286),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[25][6] ));
 DLH_X1 _12919_ (.D(net278),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[25][7] ));
 DLH_X1 _12920_ (.D(net318),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[10][0] ));
 DLH_X1 _12921_ (.D(net314),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[10][1] ));
 DLH_X1 _12922_ (.D(net309),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[10][2] ));
 DLH_X1 _12923_ (.D(net301),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[10][3] ));
 DLH_X1 _12924_ (.D(net296),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[10][4] ));
 DLH_X1 _12925_ (.D(net290),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[10][5] ));
 DLH_X1 _12926_ (.D(net286),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[10][6] ));
 DLH_X1 _12927_ (.D(net278),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[10][7] ));
 DLH_X1 _12928_ (.D(net319),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[3][0] ));
 DLH_X1 _12929_ (.D(net314),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[3][1] ));
 DLH_X1 _12930_ (.D(net309),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[3][2] ));
 DLH_X1 _12931_ (.D(net301),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[3][3] ));
 DLH_X1 _12932_ (.D(net296),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[3][4] ));
 DLH_X1 _12933_ (.D(net290),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[3][5] ));
 DLH_X1 _12934_ (.D(net286),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[3][6] ));
 DLH_X1 _12935_ (.D(net279),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[3][7] ));
 DLH_X1 _12936_ (.D(net319),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[16][0] ));
 DLH_X1 _12937_ (.D(net314),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[16][1] ));
 DLH_X1 _12938_ (.D(net307),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[16][2] ));
 DLH_X1 _12939_ (.D(net301),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[16][3] ));
 DLH_X1 _12940_ (.D(net296),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[16][4] ));
 DLH_X1 _12941_ (.D(net290),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[16][5] ));
 DLH_X1 _12942_ (.D(net286),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[16][6] ));
 DLH_X1 _12943_ (.D(net278),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[16][7] ));
 DLH_X1 _12944_ (.D(net319),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[24][0] ));
 DLH_X1 _12945_ (.D(net314),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[24][1] ));
 DLH_X1 _12946_ (.D(net307),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[24][2] ));
 DLH_X1 _12947_ (.D(net301),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[24][3] ));
 DLH_X1 _12948_ (.D(net296),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[24][4] ));
 DLH_X1 _12949_ (.D(net290),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[24][5] ));
 DLH_X1 _12950_ (.D(net286),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[24][6] ));
 DLH_X1 _12951_ (.D(net279),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[24][7] ));
 DLH_X1 _12952_ (.D(net318),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[4][0] ));
 DLH_X1 _12953_ (.D(net314),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[4][1] ));
 DLH_X1 _12954_ (.D(net307),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[4][2] ));
 DLH_X1 _12955_ (.D(net301),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[4][3] ));
 DLH_X1 _12956_ (.D(net296),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[4][4] ));
 DLH_X1 _12957_ (.D(net290),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[4][5] ));
 DLH_X1 _12958_ (.D(net281),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[4][6] ));
 DLH_X1 _12959_ (.D(net278),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[4][7] ));
 DLH_X1 _12960_ (.D(net319),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[15][0] ));
 DLH_X1 _12961_ (.D(net314),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[15][1] ));
 DLH_X1 _12962_ (.D(net307),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[15][2] ));
 DLH_X1 _12963_ (.D(net301),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[15][3] ));
 DLH_X1 _12964_ (.D(net296),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[15][4] ));
 DLH_X1 _12965_ (.D(net290),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[15][5] ));
 DLH_X1 _12966_ (.D(net286),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[15][6] ));
 DLH_X1 _12967_ (.D(net279),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[15][7] ));
 DLH_X1 _12968_ (.D(net318),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[11][0] ));
 DLH_X1 _12969_ (.D(net313),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[11][1] ));
 DLH_X1 _12970_ (.D(net309),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[11][2] ));
 DLH_X1 _12971_ (.D(net301),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[11][3] ));
 DLH_X1 _12972_ (.D(net296),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[11][4] ));
 DLH_X1 _12973_ (.D(net290),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[11][5] ));
 DLH_X1 _12974_ (.D(net286),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[11][6] ));
 DLH_X1 _12975_ (.D(net278),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[11][7] ));
 DLH_X1 _12976_ (.D(net319),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[5][0] ));
 DLH_X1 _12977_ (.D(net314),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[5][1] ));
 DLH_X1 _12978_ (.D(net307),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[5][2] ));
 DLH_X1 _12979_ (.D(net301),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[5][3] ));
 DLH_X1 _12980_ (.D(net296),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[5][4] ));
 DLH_X1 _12981_ (.D(net290),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[5][5] ));
 DLH_X1 _12982_ (.D(net286),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[5][6] ));
 DLH_X1 _12983_ (.D(net278),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[5][7] ));
 DLH_X1 _12984_ (.D(net319),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[23][0] ));
 DLH_X1 _12985_ (.D(net314),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[23][1] ));
 DLH_X1 _12986_ (.D(net307),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[23][2] ));
 DLH_X1 _12987_ (.D(net301),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[23][3] ));
 DLH_X1 _12988_ (.D(net296),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[23][4] ));
 DLH_X1 _12989_ (.D(net290),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[23][5] ));
 DLH_X1 _12990_ (.D(net286),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[23][6] ));
 DLH_X1 _12991_ (.D(net279),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[23][7] ));
 DLH_X1 _12992_ (.D(net319),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[19][0] ));
 DLH_X1 _12993_ (.D(net314),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[19][1] ));
 DLH_X1 _12994_ (.D(net309),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[19][2] ));
 DLH_X1 _12995_ (.D(net301),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[19][3] ));
 DLH_X1 _12996_ (.D(net296),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[19][4] ));
 DLH_X1 _12997_ (.D(net290),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[19][5] ));
 DLH_X1 _12998_ (.D(net281),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[19][6] ));
 DLH_X1 _12999_ (.D(net279),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[19][7] ));
 DLH_X1 _13000_ (.D(net319),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[31][0] ));
 DLH_X1 _13001_ (.D(net314),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[31][1] ));
 DLH_X1 _13002_ (.D(net309),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[31][2] ));
 DLH_X1 _13003_ (.D(net301),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[31][3] ));
 DLH_X1 _13004_ (.D(net296),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[31][4] ));
 DLH_X1 _13005_ (.D(net290),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[31][5] ));
 DLH_X1 _13006_ (.D(net281),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[31][6] ));
 DLH_X1 _13007_ (.D(net278),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[31][7] ));
 DLH_X1 _13008_ (.D(net319),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[6][0] ));
 DLH_X1 _13009_ (.D(net314),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[6][1] ));
 DLH_X1 _13010_ (.D(net309),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[6][2] ));
 DLH_X1 _13011_ (.D(net301),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[6][3] ));
 DLH_X1 _13012_ (.D(net296),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[6][4] ));
 DLH_X1 _13013_ (.D(net289),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[6][5] ));
 DLH_X1 _13014_ (.D(net286),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[6][6] ));
 DLH_X1 _13015_ (.D(net278),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[6][7] ));
 DLH_X1 _13016_ (.D(net318),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[14][0] ));
 DLH_X1 _13017_ (.D(net313),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[14][1] ));
 DLH_X1 _13018_ (.D(net307),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[14][2] ));
 DLH_X1 _13019_ (.D(net301),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[14][3] ));
 DLH_X1 _13020_ (.D(net296),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[14][4] ));
 DLH_X1 _13021_ (.D(net290),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[14][5] ));
 DLH_X1 _13022_ (.D(net286),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[14][6] ));
 DLH_X1 _13023_ (.D(net278),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[14][7] ));
 DLH_X1 _13024_ (.D(net318),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[30][0] ));
 DLH_X1 _13025_ (.D(net314),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[30][1] ));
 DLH_X1 _13026_ (.D(net307),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[30][2] ));
 DLH_X1 _13027_ (.D(net301),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[30][3] ));
 DLH_X1 _13028_ (.D(net296),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[30][4] ));
 DLH_X1 _13029_ (.D(net290),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[30][5] ));
 DLH_X1 _13030_ (.D(net286),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[30][6] ));
 DLH_X1 _13031_ (.D(net279),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[30][7] ));
 DLH_X1 _13032_ (.D(net319),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[22][0] ));
 DLH_X1 _13033_ (.D(net314),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[22][1] ));
 DLH_X1 _13034_ (.D(net307),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[22][2] ));
 DLH_X1 _13035_ (.D(net301),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[22][3] ));
 DLH_X1 _13036_ (.D(net296),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[22][4] ));
 DLH_X1 _13037_ (.D(net290),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[22][5] ));
 DLH_X1 _13038_ (.D(net286),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[22][6] ));
 DLH_X1 _13039_ (.D(net279),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[22][7] ));
 DLH_X1 _13040_ (.D(net318),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[7][0] ));
 DLH_X1 _13041_ (.D(net314),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[7][1] ));
 DLH_X1 _13042_ (.D(net309),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[7][2] ));
 DLH_X1 _13043_ (.D(net301),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[7][3] ));
 DLH_X1 _13044_ (.D(net296),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[7][4] ));
 DLH_X1 _13045_ (.D(net290),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[7][5] ));
 DLH_X1 _13046_ (.D(net286),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[7][6] ));
 DLH_X1 _13047_ (.D(net279),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[7][7] ));
 DLH_X1 _13048_ (.D(net318),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[29][0] ));
 DLH_X1 _13049_ (.D(net313),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[29][1] ));
 DLH_X1 _13050_ (.D(net307),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[29][2] ));
 DLH_X1 _13051_ (.D(net301),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[29][3] ));
 DLH_X1 _13052_ (.D(net296),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[29][4] ));
 DLH_X1 _13053_ (.D(net290),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[29][5] ));
 DLH_X1 _13054_ (.D(net286),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[29][6] ));
 DLH_X1 _13055_ (.D(net279),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[29][7] ));
 DLH_X1 _13056_ (.D(net318),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[12][0] ));
 DLH_X1 _13057_ (.D(net314),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[12][1] ));
 DLH_X1 _13058_ (.D(net307),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[12][2] ));
 DLH_X1 _13059_ (.D(net301),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[12][3] ));
 DLH_X1 _13060_ (.D(net296),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[12][4] ));
 DLH_X1 _13061_ (.D(net289),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[12][5] ));
 DLH_X1 _13062_ (.D(net286),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[12][6] ));
 DLH_X1 _13063_ (.D(net279),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[12][7] ));
 DLH_X1 _13064_ (.D(net319),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[17][0] ));
 DLH_X1 _13065_ (.D(net314),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[17][1] ));
 DLH_X1 _13066_ (.D(net309),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[17][2] ));
 DLH_X1 _13067_ (.D(net301),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[17][3] ));
 DLH_X1 _13068_ (.D(net296),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[17][4] ));
 DLH_X1 _13069_ (.D(net290),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[17][5] ));
 DLH_X1 _13070_ (.D(net286),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[17][6] ));
 DLH_X1 _13071_ (.D(net279),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[17][7] ));
 DLH_X1 _13072_ (.D(net319),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[28][0] ));
 DLH_X1 _13073_ (.D(net314),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[28][1] ));
 DLH_X1 _13074_ (.D(net309),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[28][2] ));
 DLH_X1 _13075_ (.D(net301),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[28][3] ));
 DLH_X1 _13076_ (.D(net296),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[28][4] ));
 DLH_X1 _13077_ (.D(net290),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[28][5] ));
 DLH_X1 _13078_ (.D(net286),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[28][6] ));
 DLH_X1 _13079_ (.D(net279),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[28][7] ));
 DLH_X1 _13080_ (.D(net318),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[8][0] ));
 DLH_X1 _13081_ (.D(net314),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[8][1] ));
 DLH_X1 _13082_ (.D(net307),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[8][2] ));
 DLH_X1 _13083_ (.D(net301),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[8][3] ));
 DLH_X1 _13084_ (.D(net296),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[8][4] ));
 DLH_X1 _13085_ (.D(net289),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[8][5] ));
 DLH_X1 _13086_ (.D(net286),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[8][6] ));
 DLH_X1 _13087_ (.D(net278),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[8][7] ));
 DLH_X1 _13088_ (.D(net319),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[21][0] ));
 DLH_X1 _13089_ (.D(net313),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[21][1] ));
 DLH_X1 _13090_ (.D(net307),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[21][2] ));
 DLH_X1 _13091_ (.D(net301),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[21][3] ));
 DLH_X1 _13092_ (.D(net296),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[21][4] ));
 DLH_X1 _13093_ (.D(net290),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[21][5] ));
 DLH_X1 _13094_ (.D(net286),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[21][6] ));
 DLH_X1 _13095_ (.D(net278),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[21][7] ));
 DLH_X1 _13096_ (.D(net319),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[27][0] ));
 DLH_X1 _13097_ (.D(net314),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[27][1] ));
 DLH_X1 _13098_ (.D(net309),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[27][2] ));
 DLH_X1 _13099_ (.D(net301),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[27][3] ));
 DLH_X1 _13100_ (.D(net296),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[27][4] ));
 DLH_X1 _13101_ (.D(net289),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[27][5] ));
 DLH_X1 _13102_ (.D(net286),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[27][6] ));
 DLH_X1 _13103_ (.D(net278),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[27][7] ));
 DLH_X1 _13104_ (.D(net318),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[18][0] ));
 DLH_X1 _13105_ (.D(net314),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[18][1] ));
 DLH_X1 _13106_ (.D(net309),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[18][2] ));
 DLH_X1 _13107_ (.D(net301),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[18][3] ));
 DLH_X1 _13108_ (.D(net296),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[18][4] ));
 DLH_X1 _13109_ (.D(net290),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[18][5] ));
 DLH_X1 _13110_ (.D(net286),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[18][6] ));
 DLH_X1 _13111_ (.D(net278),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.mem[18][7] ));
 DLL_X1 _13112_ (.D(\lut.gen_sub_units_scm.__4.sub_unit_i.cg_we_global.en_i ),
    .GN(clknet_level_5_1_2116__00532_),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.cg_we_global.clk_en ));
 DLL_X1 _13113_ (.D(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__0.cg_i.en_i ),
    .GN(clknet_level_2_1_5203__00567_),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_en ));
 DLL_X1 _13114_ (.D(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__1.cg_i.en_i ),
    .GN(clknet_level_2_1_4200__00567_),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_en ));
 DLL_X1 _13115_ (.D(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__2.cg_i.en_i ),
    .GN(clknet_level_2_1_1191__00567_),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_en ));
 DLL_X1 _13116_ (.D(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__3.cg_i.en_i ),
    .GN(clknet_level_2_1_7209__00567_),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_en ));
 DLL_X1 _13117_ (.D(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__4.cg_i.en_i ),
    .GN(clknet_level_2_1_3197__00567_),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_en ));
 DLL_X1 _13118_ (.D(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__5.cg_i.en_i ),
    .GN(clknet_level_2_1_4200__00567_),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_en ));
 DLL_X1 _13119_ (.D(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__6.cg_i.en_i ),
    .GN(clknet_level_2_1_8212__00567_),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_en ));
 DLL_X1 _13120_ (.D(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__7.cg_i.en_i ),
    .GN(clknet_level_2_1_6206__00567_),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_en ));
 DLL_X1 _13121_ (.D(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__8.cg_i.en_i ),
    .GN(clknet_level_2_1_3197__00567_),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_en ));
 DLL_X1 _13122_ (.D(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__9.cg_i.en_i ),
    .GN(clknet_level_2_1_3197__00567_),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_en ));
 DLL_X1 _13123_ (.D(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__10.cg_i.en_i ),
    .GN(clknet_level_2_1_1191__00567_),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_en ));
 DLL_X1 _13124_ (.D(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__11.cg_i.en_i ),
    .GN(clknet_level_2_1_3197__00567_),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_en ));
 DLL_X1 _13125_ (.D(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__12.cg_i.en_i ),
    .GN(clknet_level_2_1_1191__00567_),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_en ));
 DLL_X1 _13126_ (.D(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__13.cg_i.en_i ),
    .GN(clknet_level_2_1_7209__00567_),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_en ));
 DLL_X1 _13127_ (.D(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__14.cg_i.en_i ),
    .GN(clknet_level_2_1_2194__00567_),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_en ));
 DLL_X1 _13128_ (.D(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__15.cg_i.en_i ),
    .GN(clknet_level_2_1_6206__00567_),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_en ));
 DLL_X1 _13129_ (.D(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__16.cg_i.en_i ),
    .GN(clknet_level_2_1_7209__00567_),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_en ));
 DLL_X1 _13130_ (.D(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__17.cg_i.en_i ),
    .GN(clknet_level_2_1_8212__00567_),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_en ));
 DLL_X1 _13131_ (.D(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__18.cg_i.en_i ),
    .GN(clknet_level_2_1_7209__00567_),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_en ));
 DLL_X1 _13132_ (.D(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__19.cg_i.en_i ),
    .GN(clknet_level_2_1_7209__00567_),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_en ));
 DLL_X1 _13133_ (.D(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__20.cg_i.en_i ),
    .GN(clknet_level_2_1_8212__00567_),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_en ));
 DLL_X1 _13134_ (.D(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__21.cg_i.en_i ),
    .GN(clknet_level_2_1_4200__00567_),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_en ));
 DLL_X1 _13135_ (.D(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__22.cg_i.en_i ),
    .GN(clknet_level_2_1_6206__00567_),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_en ));
 DLL_X1 _13136_ (.D(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__23.cg_i.en_i ),
    .GN(clknet_level_2_1_8212__00567_),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_en ));
 DLL_X1 _13137_ (.D(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__24.cg_i.en_i ),
    .GN(clknet_level_2_1_4200__00567_),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_en ));
 DLL_X1 _13138_ (.D(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__25.cg_i.en_i ),
    .GN(clknet_level_2_1_4200__00567_),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_en ));
 DLL_X1 _13139_ (.D(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__26.cg_i.en_i ),
    .GN(clknet_level_2_1_1191__00567_),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_en ));
 DLL_X1 _13140_ (.D(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__27.cg_i.en_i ),
    .GN(clknet_level_2_1_4200__00567_),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_en ));
 DLL_X1 _13141_ (.D(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__28.cg_i.en_i ),
    .GN(clknet_level_2_1_8212__00567_),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_en ));
 DLL_X1 _13142_ (.D(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__29.cg_i.en_i ),
    .GN(clknet_level_2_1_5203__00567_),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_en ));
 DLL_X1 _13143_ (.D(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__30.cg_i.en_i ),
    .GN(clknet_level_2_1_5203__00567_),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_en ));
 DLL_X1 _13144_ (.D(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__31.cg_i.en_i ),
    .GN(clknet_level_2_1_3197__00567_),
    .Q(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_en ));
 DLH_X1 _13145_ (.D(net317),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[13][0] ));
 DLH_X1 _13146_ (.D(net311),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[13][1] ));
 DLH_X1 _13147_ (.D(net305),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[13][2] ));
 DLH_X1 _13148_ (.D(net299),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[13][3] ));
 DLH_X1 _13149_ (.D(net293),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[13][4] ));
 DLH_X1 _13150_ (.D(net287),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[13][5] ));
 DLH_X1 _13151_ (.D(net284),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[13][6] ));
 DLH_X1 _13152_ (.D(net275),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[13][7] ));
 DLH_X1 _13153_ (.D(net320),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[1][0] ));
 DLH_X1 _13154_ (.D(net311),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[1][1] ));
 DLH_X1 _13155_ (.D(net305),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[1][2] ));
 DLH_X1 _13156_ (.D(net299),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[1][3] ));
 DLH_X1 _13157_ (.D(net293),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[1][4] ));
 DLH_X1 _13158_ (.D(net287),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[1][5] ));
 DLH_X1 _13159_ (.D(net284),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[1][6] ));
 DLH_X1 _13160_ (.D(net275),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[1][7] ));
 DLH_X1 _13161_ (.D(net317),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[26][0] ));
 DLH_X1 _13162_ (.D(net311),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[26][1] ));
 DLH_X1 _13163_ (.D(net305),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[26][2] ));
 DLH_X1 _13164_ (.D(net299),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[26][3] ));
 DLH_X1 _13165_ (.D(net293),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[26][4] ));
 DLH_X1 _13166_ (.D(net287),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[26][5] ));
 DLH_X1 _13167_ (.D(net284),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[26][6] ));
 DLH_X1 _13168_ (.D(net275),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[26][7] ));
 DLH_X1 _13169_ (.D(net317),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[9][0] ));
 DLH_X1 _13170_ (.D(net310),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[9][1] ));
 DLH_X1 _13171_ (.D(net305),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[9][2] ));
 DLH_X1 _13172_ (.D(net299),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[9][3] ));
 DLH_X1 _13173_ (.D(net293),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[9][4] ));
 DLH_X1 _13174_ (.D(net287),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[9][5] ));
 DLH_X1 _13175_ (.D(net284),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[9][6] ));
 DLH_X1 _13176_ (.D(net275),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[9][7] ));
 DLH_X1 _13177_ (.D(net317),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[0][0] ));
 DLH_X1 _13178_ (.D(net311),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[0][1] ));
 DLH_X1 _13179_ (.D(net306),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[0][2] ));
 DLH_X1 _13180_ (.D(net303),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[0][3] ));
 DLH_X1 _13181_ (.D(net294),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[0][4] ));
 DLH_X1 _13182_ (.D(net292),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[0][5] ));
 DLH_X1 _13183_ (.D(net284),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[0][6] ));
 DLH_X1 _13184_ (.D(net277),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[0][7] ));
 DLH_X1 _13185_ (.D(net317),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[20][0] ));
 DLH_X1 _13186_ (.D(net311),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[20][1] ));
 DLH_X1 _13187_ (.D(net305),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[20][2] ));
 DLH_X1 _13188_ (.D(net299),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[20][3] ));
 DLH_X1 _13189_ (.D(net293),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[20][4] ));
 DLH_X1 _13190_ (.D(net287),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[20][5] ));
 DLH_X1 _13191_ (.D(net284),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[20][6] ));
 DLH_X1 _13192_ (.D(net275),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[20][7] ));
 DLH_X1 _13193_ (.D(net320),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[2][0] ));
 DLH_X1 _13194_ (.D(net310),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[2][1] ));
 DLH_X1 _13195_ (.D(net305),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[2][2] ));
 DLH_X1 _13196_ (.D(net299),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[2][3] ));
 DLH_X1 _13197_ (.D(net293),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[2][4] ));
 DLH_X1 _13198_ (.D(net287),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[2][5] ));
 DLH_X1 _13199_ (.D(net284),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[2][6] ));
 DLH_X1 _13200_ (.D(net275),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[2][7] ));
 DLH_X1 _13201_ (.D(net317),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[25][0] ));
 DLH_X1 _13202_ (.D(net311),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[25][1] ));
 DLH_X1 _13203_ (.D(net305),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[25][2] ));
 DLH_X1 _13204_ (.D(net299),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[25][3] ));
 DLH_X1 _13205_ (.D(net293),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[25][4] ));
 DLH_X1 _13206_ (.D(net287),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[25][5] ));
 DLH_X1 _13207_ (.D(net284),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[25][6] ));
 DLH_X1 _13208_ (.D(net275),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[25][7] ));
 DLH_X1 _13209_ (.D(net320),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[10][0] ));
 DLH_X1 _13210_ (.D(net310),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[10][1] ));
 DLH_X1 _13211_ (.D(net305),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[10][2] ));
 DLH_X1 _13212_ (.D(net299),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[10][3] ));
 DLH_X1 _13213_ (.D(net293),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[10][4] ));
 DLH_X1 _13214_ (.D(net287),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[10][5] ));
 DLH_X1 _13215_ (.D(net284),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[10][6] ));
 DLH_X1 _13216_ (.D(net275),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[10][7] ));
 DLH_X1 _13217_ (.D(net320),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[3][0] ));
 DLH_X1 _13218_ (.D(net311),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[3][1] ));
 DLH_X1 _13219_ (.D(net305),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[3][2] ));
 DLH_X1 _13220_ (.D(net299),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[3][3] ));
 DLH_X1 _13221_ (.D(net293),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[3][4] ));
 DLH_X1 _13222_ (.D(net287),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[3][5] ));
 DLH_X1 _13223_ (.D(net284),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[3][6] ));
 DLH_X1 _13224_ (.D(net275),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[3][7] ));
 DLH_X1 _13225_ (.D(net317),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[16][0] ));
 DLH_X1 _13226_ (.D(net311),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[16][1] ));
 DLH_X1 _13227_ (.D(net305),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[16][2] ));
 DLH_X1 _13228_ (.D(net299),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[16][3] ));
 DLH_X1 _13229_ (.D(net293),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[16][4] ));
 DLH_X1 _13230_ (.D(net287),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[16][5] ));
 DLH_X1 _13231_ (.D(net284),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[16][6] ));
 DLH_X1 _13232_ (.D(net275),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[16][7] ));
 DLH_X1 _13233_ (.D(net317),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[24][0] ));
 DLH_X1 _13234_ (.D(net311),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[24][1] ));
 DLH_X1 _13235_ (.D(net305),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[24][2] ));
 DLH_X1 _13236_ (.D(net299),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[24][3] ));
 DLH_X1 _13237_ (.D(net293),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[24][4] ));
 DLH_X1 _13238_ (.D(net287),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[24][5] ));
 DLH_X1 _13239_ (.D(net284),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[24][6] ));
 DLH_X1 _13240_ (.D(net275),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[24][7] ));
 DLH_X1 _13241_ (.D(net320),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[4][0] ));
 DLH_X1 _13242_ (.D(net311),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[4][1] ));
 DLH_X1 _13243_ (.D(net305),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[4][2] ));
 DLH_X1 _13244_ (.D(net299),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[4][3] ));
 DLH_X1 _13245_ (.D(net293),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[4][4] ));
 DLH_X1 _13246_ (.D(net287),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[4][5] ));
 DLH_X1 _13247_ (.D(net284),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[4][6] ));
 DLH_X1 _13248_ (.D(net275),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[4][7] ));
 DLH_X1 _13249_ (.D(net320),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[15][0] ));
 DLH_X1 _13250_ (.D(net311),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[15][1] ));
 DLH_X1 _13251_ (.D(net305),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[15][2] ));
 DLH_X1 _13252_ (.D(net299),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[15][3] ));
 DLH_X1 _13253_ (.D(net293),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[15][4] ));
 DLH_X1 _13254_ (.D(net287),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[15][5] ));
 DLH_X1 _13255_ (.D(net284),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[15][6] ));
 DLH_X1 _13256_ (.D(net275),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[15][7] ));
 DLH_X1 _13257_ (.D(net320),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[11][0] ));
 DLH_X1 _13258_ (.D(net311),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[11][1] ));
 DLH_X1 _13259_ (.D(net305),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[11][2] ));
 DLH_X1 _13260_ (.D(net299),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[11][3] ));
 DLH_X1 _13261_ (.D(net293),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[11][4] ));
 DLH_X1 _13262_ (.D(net287),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[11][5] ));
 DLH_X1 _13263_ (.D(net284),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[11][6] ));
 DLH_X1 _13264_ (.D(net275),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[11][7] ));
 DLH_X1 _13265_ (.D(net317),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[5][0] ));
 DLH_X1 _13266_ (.D(net311),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[5][1] ));
 DLH_X1 _13267_ (.D(net305),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[5][2] ));
 DLH_X1 _13268_ (.D(net299),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[5][3] ));
 DLH_X1 _13269_ (.D(net293),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[5][4] ));
 DLH_X1 _13270_ (.D(net287),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[5][5] ));
 DLH_X1 _13271_ (.D(net284),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[5][6] ));
 DLH_X1 _13272_ (.D(net275),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[5][7] ));
 DLH_X1 _13273_ (.D(net317),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[23][0] ));
 DLH_X1 _13274_ (.D(net311),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[23][1] ));
 DLH_X1 _13275_ (.D(net305),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[23][2] ));
 DLH_X1 _13276_ (.D(net299),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[23][3] ));
 DLH_X1 _13277_ (.D(net293),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[23][4] ));
 DLH_X1 _13278_ (.D(net287),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[23][5] ));
 DLH_X1 _13279_ (.D(net284),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[23][6] ));
 DLH_X1 _13280_ (.D(net275),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[23][7] ));
 DLH_X1 _13281_ (.D(net320),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[19][0] ));
 DLH_X1 _13282_ (.D(net310),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[19][1] ));
 DLH_X1 _13283_ (.D(net305),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[19][2] ));
 DLH_X1 _13284_ (.D(net299),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[19][3] ));
 DLH_X1 _13285_ (.D(net293),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[19][4] ));
 DLH_X1 _13286_ (.D(net287),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[19][5] ));
 DLH_X1 _13287_ (.D(net284),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[19][6] ));
 DLH_X1 _13288_ (.D(net275),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[19][7] ));
 DLH_X1 _13289_ (.D(net320),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[31][0] ));
 DLH_X1 _13290_ (.D(net311),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[31][1] ));
 DLH_X1 _13291_ (.D(net305),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[31][2] ));
 DLH_X1 _13292_ (.D(net299),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[31][3] ));
 DLH_X1 _13293_ (.D(net293),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[31][4] ));
 DLH_X1 _13294_ (.D(net287),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[31][5] ));
 DLH_X1 _13295_ (.D(net284),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[31][6] ));
 DLH_X1 _13296_ (.D(net275),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[31][7] ));
 DLH_X1 _13297_ (.D(net317),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[6][0] ));
 DLH_X1 _13298_ (.D(net311),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[6][1] ));
 DLH_X1 _13299_ (.D(net305),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[6][2] ));
 DLH_X1 _13300_ (.D(net299),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[6][3] ));
 DLH_X1 _13301_ (.D(net293),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[6][4] ));
 DLH_X1 _13302_ (.D(net287),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[6][5] ));
 DLH_X1 _13303_ (.D(net284),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[6][6] ));
 DLH_X1 _13304_ (.D(net275),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[6][7] ));
 DLH_X1 _13305_ (.D(net320),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[14][0] ));
 DLH_X1 _13306_ (.D(net311),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[14][1] ));
 DLH_X1 _13307_ (.D(net305),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[14][2] ));
 DLH_X1 _13308_ (.D(net299),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[14][3] ));
 DLH_X1 _13309_ (.D(net293),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[14][4] ));
 DLH_X1 _13310_ (.D(net287),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[14][5] ));
 DLH_X1 _13311_ (.D(net284),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[14][6] ));
 DLH_X1 _13312_ (.D(net275),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[14][7] ));
 DLH_X1 _13313_ (.D(net320),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[30][0] ));
 DLH_X1 _13314_ (.D(net311),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[30][1] ));
 DLH_X1 _13315_ (.D(net305),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[30][2] ));
 DLH_X1 _13316_ (.D(net299),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[30][3] ));
 DLH_X1 _13317_ (.D(net293),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[30][4] ));
 DLH_X1 _13318_ (.D(net287),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[30][5] ));
 DLH_X1 _13319_ (.D(net284),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[30][6] ));
 DLH_X1 _13320_ (.D(net275),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[30][7] ));
 DLH_X1 _13321_ (.D(net320),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[22][0] ));
 DLH_X1 _13322_ (.D(net311),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[22][1] ));
 DLH_X1 _13323_ (.D(net305),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[22][2] ));
 DLH_X1 _13324_ (.D(net299),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[22][3] ));
 DLH_X1 _13325_ (.D(net293),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[22][4] ));
 DLH_X1 _13326_ (.D(net287),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[22][5] ));
 DLH_X1 _13327_ (.D(net284),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[22][6] ));
 DLH_X1 _13328_ (.D(net275),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[22][7] ));
 DLH_X1 _13329_ (.D(net317),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[7][0] ));
 DLH_X1 _13330_ (.D(net311),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[7][1] ));
 DLH_X1 _13331_ (.D(net305),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[7][2] ));
 DLH_X1 _13332_ (.D(net299),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[7][3] ));
 DLH_X1 _13333_ (.D(net293),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[7][4] ));
 DLH_X1 _13334_ (.D(net287),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[7][5] ));
 DLH_X1 _13335_ (.D(net284),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[7][6] ));
 DLH_X1 _13336_ (.D(net275),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[7][7] ));
 DLH_X1 _13337_ (.D(net320),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[29][0] ));
 DLH_X1 _13338_ (.D(net311),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[29][1] ));
 DLH_X1 _13339_ (.D(net305),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[29][2] ));
 DLH_X1 _13340_ (.D(net299),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[29][3] ));
 DLH_X1 _13341_ (.D(net293),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[29][4] ));
 DLH_X1 _13342_ (.D(net287),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[29][5] ));
 DLH_X1 _13343_ (.D(net284),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[29][6] ));
 DLH_X1 _13344_ (.D(net275),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[29][7] ));
 DLH_X1 _13345_ (.D(net317),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[12][0] ));
 DLH_X1 _13346_ (.D(net311),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[12][1] ));
 DLH_X1 _13347_ (.D(net305),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[12][2] ));
 DLH_X1 _13348_ (.D(net299),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[12][3] ));
 DLH_X1 _13349_ (.D(net293),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[12][4] ));
 DLH_X1 _13350_ (.D(net287),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[12][5] ));
 DLH_X1 _13351_ (.D(net284),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[12][6] ));
 DLH_X1 _13352_ (.D(net275),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[12][7] ));
 DLH_X1 _13353_ (.D(net317),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[17][0] ));
 DLH_X1 _13354_ (.D(net310),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[17][1] ));
 DLH_X1 _13355_ (.D(net305),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[17][2] ));
 DLH_X1 _13356_ (.D(net299),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[17][3] ));
 DLH_X1 _13357_ (.D(net293),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[17][4] ));
 DLH_X1 _13358_ (.D(net287),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[17][5] ));
 DLH_X1 _13359_ (.D(net284),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[17][6] ));
 DLH_X1 _13360_ (.D(net275),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[17][7] ));
 DLH_X1 _13361_ (.D(net317),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[28][0] ));
 DLH_X1 _13362_ (.D(net311),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[28][1] ));
 DLH_X1 _13363_ (.D(net305),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[28][2] ));
 DLH_X1 _13364_ (.D(net299),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[28][3] ));
 DLH_X1 _13365_ (.D(net293),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[28][4] ));
 DLH_X1 _13366_ (.D(net287),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[28][5] ));
 DLH_X1 _13367_ (.D(net284),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[28][6] ));
 DLH_X1 _13368_ (.D(net275),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[28][7] ));
 DLH_X1 _13369_ (.D(net320),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[8][0] ));
 DLH_X1 _13370_ (.D(net310),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[8][1] ));
 DLH_X1 _13371_ (.D(net305),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[8][2] ));
 DLH_X1 _13372_ (.D(net299),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[8][3] ));
 DLH_X1 _13373_ (.D(net293),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[8][4] ));
 DLH_X1 _13374_ (.D(net287),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[8][5] ));
 DLH_X1 _13375_ (.D(net284),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[8][6] ));
 DLH_X1 _13376_ (.D(net275),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[8][7] ));
 DLH_X1 _13377_ (.D(net317),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[21][0] ));
 DLH_X1 _13378_ (.D(net311),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[21][1] ));
 DLH_X1 _13379_ (.D(net305),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[21][2] ));
 DLH_X1 _13380_ (.D(net299),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[21][3] ));
 DLH_X1 _13381_ (.D(net293),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[21][4] ));
 DLH_X1 _13382_ (.D(net287),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[21][5] ));
 DLH_X1 _13383_ (.D(net284),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[21][6] ));
 DLH_X1 _13384_ (.D(net275),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[21][7] ));
 DLH_X1 _13385_ (.D(net320),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[27][0] ));
 DLH_X1 _13386_ (.D(net310),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[27][1] ));
 DLH_X1 _13387_ (.D(net305),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[27][2] ));
 DLH_X1 _13388_ (.D(net299),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[27][3] ));
 DLH_X1 _13389_ (.D(net293),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[27][4] ));
 DLH_X1 _13390_ (.D(net287),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[27][5] ));
 DLH_X1 _13391_ (.D(net284),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[27][6] ));
 DLH_X1 _13392_ (.D(net275),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[27][7] ));
 DLH_X1 _13393_ (.D(net320),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[18][0] ));
 DLH_X1 _13394_ (.D(net310),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[18][1] ));
 DLH_X1 _13395_ (.D(net305),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[18][2] ));
 DLH_X1 _13396_ (.D(net299),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[18][3] ));
 DLH_X1 _13397_ (.D(net293),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[18][4] ));
 DLH_X1 _13398_ (.D(net287),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[18][5] ));
 DLH_X1 _13399_ (.D(net284),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[18][6] ));
 DLH_X1 _13400_ (.D(net275),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.mem[18][7] ));
 DLL_X1 _13401_ (.D(\lut.gen_sub_units_scm.__3.sub_unit_i.cg_we_global.en_i ),
    .GN(clknet_level_5_1_3218__00532_),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.cg_we_global.clk_en ));
 DLL_X1 _13402_ (.D(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__0.cg_i.en_i ),
    .GN(clknet_level_2_1_8290__00570_),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_en ));
 DLL_X1 _13403_ (.D(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__1.cg_i.en_i ),
    .GN(clknet_level_2_1_2272__00570_),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_en ));
 DLL_X1 _13404_ (.D(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__2.cg_i.en_i ),
    .GN(clknet_level_2_1_4278__00570_),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_en ));
 DLL_X1 _13405_ (.D(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__3.cg_i.en_i ),
    .GN(clknet_level_2_1_2272__00570_),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_en ));
 DLL_X1 _13406_ (.D(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__4.cg_i.en_i ),
    .GN(clknet_level_2_1_1269__00570_),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_en ));
 DLL_X1 _13407_ (.D(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__5.cg_i.en_i ),
    .GN(clknet_level_2_1_6284__00570_),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_en ));
 DLL_X1 _13408_ (.D(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__6.cg_i.en_i ),
    .GN(clknet_level_2_1_7287__00570_),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_en ));
 DLL_X1 _13409_ (.D(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__7.cg_i.en_i ),
    .GN(clknet_level_2_1_8290__00570_),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_en ));
 DLL_X1 _13410_ (.D(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__8.cg_i.en_i ),
    .GN(clknet_level_2_1_7287__00570_),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_en ));
 DLL_X1 _13411_ (.D(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__9.cg_i.en_i ),
    .GN(clknet_level_2_1_7287__00570_),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_en ));
 DLL_X1 _13412_ (.D(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__10.cg_i.en_i ),
    .GN(clknet_level_2_1_8290__00570_),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_en ));
 DLL_X1 _13413_ (.D(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__11.cg_i.en_i ),
    .GN(clknet_level_2_1_7287__00570_),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_en ));
 DLL_X1 _13414_ (.D(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__12.cg_i.en_i ),
    .GN(clknet_level_2_1_4278__00570_),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_en ));
 DLL_X1 _13415_ (.D(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__13.cg_i.en_i ),
    .GN(clknet_level_2_1_1269__00570_),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_en ));
 DLL_X1 _13416_ (.D(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__14.cg_i.en_i ),
    .GN(clknet_level_2_1_1269__00570_),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_en ));
 DLL_X1 _13417_ (.D(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__15.cg_i.en_i ),
    .GN(clknet_level_2_1_1269__00570_),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_en ));
 DLL_X1 _13418_ (.D(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__16.cg_i.en_i ),
    .GN(clknet_level_2_1_2272__00570_),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_en ));
 DLL_X1 _13419_ (.D(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__17.cg_i.en_i ),
    .GN(clknet_level_2_1_2272__00570_),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_en ));
 DLL_X1 _13420_ (.D(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__18.cg_i.en_i ),
    .GN(clknet_level_2_1_3275__00570_),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_en ));
 DLL_X1 _13421_ (.D(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__19.cg_i.en_i ),
    .GN(clknet_level_2_1_3275__00570_),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_en ));
 DLL_X1 _13422_ (.D(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__20.cg_i.en_i ),
    .GN(clknet_level_2_1_5281__00570_),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_en ));
 DLL_X1 _13423_ (.D(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__21.cg_i.en_i ),
    .GN(clknet_level_2_1_5281__00570_),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_en ));
 DLL_X1 _13424_ (.D(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__22.cg_i.en_i ),
    .GN(clknet_level_2_1_1269__00570_),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_en ));
 DLL_X1 _13425_ (.D(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__23.cg_i.en_i ),
    .GN(clknet_level_2_1_5281__00570_),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_en ));
 DLL_X1 _13426_ (.D(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__24.cg_i.en_i ),
    .GN(clknet_level_2_1_5281__00570_),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_en ));
 DLL_X1 _13427_ (.D(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__25.cg_i.en_i ),
    .GN(clknet_level_2_1_7287__00570_),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_en ));
 DLL_X1 _13428_ (.D(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__26.cg_i.en_i ),
    .GN(clknet_level_2_1_2272__00570_),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_en ));
 DLL_X1 _13429_ (.D(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__27.cg_i.en_i ),
    .GN(clknet_level_2_1_8290__00570_),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_en ));
 DLL_X1 _13430_ (.D(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__28.cg_i.en_i ),
    .GN(clknet_level_2_1_5281__00570_),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_en ));
 DLL_X1 _13431_ (.D(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__29.cg_i.en_i ),
    .GN(clknet_level_2_1_7287__00570_),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_en ));
 DLL_X1 _13432_ (.D(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__30.cg_i.en_i ),
    .GN(clknet_level_2_1_4278__00570_),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_en ));
 DLL_X1 _13433_ (.D(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__31.cg_i.en_i ),
    .GN(clknet_level_2_1_8290__00570_),
    .Q(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_en ));
 DLH_X1 _13434_ (.D(net320),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[13][0] ));
 DLH_X1 _13435_ (.D(net310),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[13][1] ));
 DLH_X1 _13436_ (.D(net308),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[13][2] ));
 DLH_X1 _13437_ (.D(net299),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[13][3] ));
 DLH_X1 _13438_ (.D(net293),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[13][4] ));
 DLH_X1 _13439_ (.D(net287),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[13][5] ));
 DLH_X1 _13440_ (.D(net285),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[13][6] ));
 DLH_X1 _13441_ (.D(net275),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[13][7] ));
 DLH_X1 _13442_ (.D(net320),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[1][0] ));
 DLH_X1 _13443_ (.D(net310),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[1][1] ));
 DLH_X1 _13444_ (.D(net308),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[1][2] ));
 DLH_X1 _13445_ (.D(net300),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[1][3] ));
 DLH_X1 _13446_ (.D(net293),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[1][4] ));
 DLH_X1 _13447_ (.D(net287),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[1][5] ));
 DLH_X1 _13448_ (.D(net283),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[1][6] ));
 DLH_X1 _13449_ (.D(net275),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[1][7] ));
 DLH_X1 _13450_ (.D(net320),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[26][0] ));
 DLH_X1 _13451_ (.D(net310),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[26][1] ));
 DLH_X1 _13452_ (.D(net308),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[26][2] ));
 DLH_X1 _13453_ (.D(net300),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[26][3] ));
 DLH_X1 _13454_ (.D(net293),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[26][4] ));
 DLH_X1 _13455_ (.D(net287),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[26][5] ));
 DLH_X1 _13456_ (.D(net283),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[26][6] ));
 DLH_X1 _13457_ (.D(net275),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[26][7] ));
 DLH_X1 _13458_ (.D(net320),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[9][0] ));
 DLH_X1 _13459_ (.D(net310),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[9][1] ));
 DLH_X1 _13460_ (.D(net308),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[9][2] ));
 DLH_X1 _13461_ (.D(net299),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[9][3] ));
 DLH_X1 _13462_ (.D(net293),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[9][4] ));
 DLH_X1 _13463_ (.D(net291),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[9][5] ));
 DLH_X1 _13464_ (.D(net285),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[9][6] ));
 DLH_X1 _13465_ (.D(net275),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[9][7] ));
 DLH_X1 _13466_ (.D(net320),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[0][0] ));
 DLH_X1 _13467_ (.D(net311),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[0][1] ));
 DLH_X1 _13468_ (.D(net305),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[0][2] ));
 DLH_X1 _13469_ (.D(net300),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[0][3] ));
 DLH_X1 _13470_ (.D(net294),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[0][4] ));
 DLH_X1 _13471_ (.D(net287),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[0][5] ));
 DLH_X1 _13472_ (.D(net285),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[0][6] ));
 DLH_X1 _13473_ (.D(net275),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[0][7] ));
 DLH_X1 _13474_ (.D(net320),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[20][0] ));
 DLH_X1 _13475_ (.D(net310),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[20][1] ));
 DLH_X1 _13476_ (.D(net308),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[20][2] ));
 DLH_X1 _13477_ (.D(net299),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[20][3] ));
 DLH_X1 _13478_ (.D(net293),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[20][4] ));
 DLH_X1 _13479_ (.D(net287),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[20][5] ));
 DLH_X1 _13480_ (.D(net285),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[20][6] ));
 DLH_X1 _13481_ (.D(net275),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[20][7] ));
 DLH_X1 _13482_ (.D(net320),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[2][0] ));
 DLH_X1 _13483_ (.D(net310),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[2][1] ));
 DLH_X1 _13484_ (.D(net308),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[2][2] ));
 DLH_X1 _13485_ (.D(net299),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[2][3] ));
 DLH_X1 _13486_ (.D(net293),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[2][4] ));
 DLH_X1 _13487_ (.D(net291),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[2][5] ));
 DLH_X1 _13488_ (.D(net283),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[2][6] ));
 DLH_X1 _13489_ (.D(net275),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[2][7] ));
 DLH_X1 _13490_ (.D(net320),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[25][0] ));
 DLH_X1 _13491_ (.D(net310),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[25][1] ));
 DLH_X1 _13492_ (.D(net308),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[25][2] ));
 DLH_X1 _13493_ (.D(net299),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[25][3] ));
 DLH_X1 _13494_ (.D(net293),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[25][4] ));
 DLH_X1 _13495_ (.D(net291),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[25][5] ));
 DLH_X1 _13496_ (.D(net285),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[25][6] ));
 DLH_X1 _13497_ (.D(net275),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[25][7] ));
 DLH_X1 _13498_ (.D(net320),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[10][0] ));
 DLH_X1 _13499_ (.D(net310),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[10][1] ));
 DLH_X1 _13500_ (.D(net308),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[10][2] ));
 DLH_X1 _13501_ (.D(net300),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[10][3] ));
 DLH_X1 _13502_ (.D(net293),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[10][4] ));
 DLH_X1 _13503_ (.D(net287),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[10][5] ));
 DLH_X1 _13504_ (.D(net285),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[10][6] ));
 DLH_X1 _13505_ (.D(net275),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[10][7] ));
 DLH_X1 _13506_ (.D(net320),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[3][0] ));
 DLH_X1 _13507_ (.D(net310),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[3][1] ));
 DLH_X1 _13508_ (.D(net305),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[3][2] ));
 DLH_X1 _13509_ (.D(net299),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[3][3] ));
 DLH_X1 _13510_ (.D(net293),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[3][4] ));
 DLH_X1 _13511_ (.D(net287),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[3][5] ));
 DLH_X1 _13512_ (.D(net285),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[3][6] ));
 DLH_X1 _13513_ (.D(net275),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[3][7] ));
 DLH_X1 _13514_ (.D(net320),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[16][0] ));
 DLH_X1 _13515_ (.D(net310),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[16][1] ));
 DLH_X1 _13516_ (.D(net305),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[16][2] ));
 DLH_X1 _13517_ (.D(net299),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[16][3] ));
 DLH_X1 _13518_ (.D(net293),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[16][4] ));
 DLH_X1 _13519_ (.D(net287),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[16][5] ));
 DLH_X1 _13520_ (.D(net283),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[16][6] ));
 DLH_X1 _13521_ (.D(net275),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[16][7] ));
 DLH_X1 _13522_ (.D(net320),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[24][0] ));
 DLH_X1 _13523_ (.D(net310),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[24][1] ));
 DLH_X1 _13524_ (.D(net308),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[24][2] ));
 DLH_X1 _13525_ (.D(net300),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[24][3] ));
 DLH_X1 _13526_ (.D(net293),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[24][4] ));
 DLH_X1 _13527_ (.D(net287),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[24][5] ));
 DLH_X1 _13528_ (.D(net285),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[24][6] ));
 DLH_X1 _13529_ (.D(net275),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[24][7] ));
 DLH_X1 _13530_ (.D(net320),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[4][0] ));
 DLH_X1 _13531_ (.D(net310),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[4][1] ));
 DLH_X1 _13532_ (.D(net308),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[4][2] ));
 DLH_X1 _13533_ (.D(net299),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[4][3] ));
 DLH_X1 _13534_ (.D(net293),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[4][4] ));
 DLH_X1 _13535_ (.D(net287),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[4][5] ));
 DLH_X1 _13536_ (.D(net285),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[4][6] ));
 DLH_X1 _13537_ (.D(net275),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[4][7] ));
 DLH_X1 _13538_ (.D(net320),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[15][0] ));
 DLH_X1 _13539_ (.D(net310),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[15][1] ));
 DLH_X1 _13540_ (.D(net305),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[15][2] ));
 DLH_X1 _13541_ (.D(net299),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[15][3] ));
 DLH_X1 _13542_ (.D(net293),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[15][4] ));
 DLH_X1 _13543_ (.D(net287),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[15][5] ));
 DLH_X1 _13544_ (.D(net285),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[15][6] ));
 DLH_X1 _13545_ (.D(net275),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[15][7] ));
 DLH_X1 _13546_ (.D(net320),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[11][0] ));
 DLH_X1 _13547_ (.D(net310),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[11][1] ));
 DLH_X1 _13548_ (.D(net308),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[11][2] ));
 DLH_X1 _13549_ (.D(net299),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[11][3] ));
 DLH_X1 _13550_ (.D(net293),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[11][4] ));
 DLH_X1 _13551_ (.D(net291),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[11][5] ));
 DLH_X1 _13552_ (.D(net285),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[11][6] ));
 DLH_X1 _13553_ (.D(net275),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[11][7] ));
 DLH_X1 _13554_ (.D(net320),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[5][0] ));
 DLH_X1 _13555_ (.D(net310),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[5][1] ));
 DLH_X1 _13556_ (.D(net308),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[5][2] ));
 DLH_X1 _13557_ (.D(net300),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[5][3] ));
 DLH_X1 _13558_ (.D(net293),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[5][4] ));
 DLH_X1 _13559_ (.D(net291),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[5][5] ));
 DLH_X1 _13560_ (.D(net285),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[5][6] ));
 DLH_X1 _13561_ (.D(net275),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[5][7] ));
 DLH_X1 _13562_ (.D(net320),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[23][0] ));
 DLH_X1 _13563_ (.D(net310),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[23][1] ));
 DLH_X1 _13564_ (.D(net305),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[23][2] ));
 DLH_X1 _13565_ (.D(net299),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[23][3] ));
 DLH_X1 _13566_ (.D(net293),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[23][4] ));
 DLH_X1 _13567_ (.D(net287),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[23][5] ));
 DLH_X1 _13568_ (.D(net283),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[23][6] ));
 DLH_X1 _13569_ (.D(net275),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[23][7] ));
 DLH_X1 _13570_ (.D(net320),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[19][0] ));
 DLH_X1 _13571_ (.D(net310),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[19][1] ));
 DLH_X1 _13572_ (.D(net308),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[19][2] ));
 DLH_X1 _13573_ (.D(net299),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[19][3] ));
 DLH_X1 _13574_ (.D(net293),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[19][4] ));
 DLH_X1 _13575_ (.D(net291),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[19][5] ));
 DLH_X1 _13576_ (.D(net283),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[19][6] ));
 DLH_X1 _13577_ (.D(net275),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[19][7] ));
 DLH_X1 _13578_ (.D(net320),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[31][0] ));
 DLH_X1 _13579_ (.D(net310),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[31][1] ));
 DLH_X1 _13580_ (.D(net305),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[31][2] ));
 DLH_X1 _13581_ (.D(net300),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[31][3] ));
 DLH_X1 _13582_ (.D(net293),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[31][4] ));
 DLH_X1 _13583_ (.D(net287),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[31][5] ));
 DLH_X1 _13584_ (.D(net283),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[31][6] ));
 DLH_X1 _13585_ (.D(net275),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[31][7] ));
 DLH_X1 _13586_ (.D(net320),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[6][0] ));
 DLH_X1 _13587_ (.D(net310),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[6][1] ));
 DLH_X1 _13588_ (.D(net308),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[6][2] ));
 DLH_X1 _13589_ (.D(net299),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[6][3] ));
 DLH_X1 _13590_ (.D(net293),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[6][4] ));
 DLH_X1 _13591_ (.D(net291),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[6][5] ));
 DLH_X1 _13592_ (.D(net285),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[6][6] ));
 DLH_X1 _13593_ (.D(net275),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[6][7] ));
 DLH_X1 _13594_ (.D(net320),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[14][0] ));
 DLH_X1 _13595_ (.D(net310),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[14][1] ));
 DLH_X1 _13596_ (.D(net308),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[14][2] ));
 DLH_X1 _13597_ (.D(net300),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[14][3] ));
 DLH_X1 _13598_ (.D(net293),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[14][4] ));
 DLH_X1 _13599_ (.D(net291),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[14][5] ));
 DLH_X1 _13600_ (.D(net283),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[14][6] ));
 DLH_X1 _13601_ (.D(net275),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[14][7] ));
 DLH_X1 _13602_ (.D(net320),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[30][0] ));
 DLH_X1 _13603_ (.D(net310),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[30][1] ));
 DLH_X1 _13604_ (.D(net308),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[30][2] ));
 DLH_X1 _13605_ (.D(net300),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[30][3] ));
 DLH_X1 _13606_ (.D(net293),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[30][4] ));
 DLH_X1 _13607_ (.D(net291),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[30][5] ));
 DLH_X1 _13608_ (.D(net285),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[30][6] ));
 DLH_X1 _13609_ (.D(net275),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[30][7] ));
 DLH_X1 _13610_ (.D(net320),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[22][0] ));
 DLH_X1 _13611_ (.D(net310),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[22][1] ));
 DLH_X1 _13612_ (.D(net308),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[22][2] ));
 DLH_X1 _13613_ (.D(net299),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[22][3] ));
 DLH_X1 _13614_ (.D(net293),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[22][4] ));
 DLH_X1 _13615_ (.D(net287),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[22][5] ));
 DLH_X1 _13616_ (.D(net283),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[22][6] ));
 DLH_X1 _13617_ (.D(net275),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[22][7] ));
 DLH_X1 _13618_ (.D(net320),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[7][0] ));
 DLH_X1 _13619_ (.D(net310),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[7][1] ));
 DLH_X1 _13620_ (.D(net305),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[7][2] ));
 DLH_X1 _13621_ (.D(net299),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[7][3] ));
 DLH_X1 _13622_ (.D(net293),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[7][4] ));
 DLH_X1 _13623_ (.D(net287),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[7][5] ));
 DLH_X1 _13624_ (.D(net283),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[7][6] ));
 DLH_X1 _13625_ (.D(net275),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[7][7] ));
 DLH_X1 _13626_ (.D(net320),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[29][0] ));
 DLH_X1 _13627_ (.D(net310),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[29][1] ));
 DLH_X1 _13628_ (.D(net308),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[29][2] ));
 DLH_X1 _13629_ (.D(net300),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[29][3] ));
 DLH_X1 _13630_ (.D(net293),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[29][4] ));
 DLH_X1 _13631_ (.D(net287),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[29][5] ));
 DLH_X1 _13632_ (.D(net283),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[29][6] ));
 DLH_X1 _13633_ (.D(net275),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[29][7] ));
 DLH_X1 _13634_ (.D(net320),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[12][0] ));
 DLH_X1 _13635_ (.D(net310),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[12][1] ));
 DLH_X1 _13636_ (.D(net308),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[12][2] ));
 DLH_X1 _13637_ (.D(net300),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[12][3] ));
 DLH_X1 _13638_ (.D(net293),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[12][4] ));
 DLH_X1 _13639_ (.D(net291),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[12][5] ));
 DLH_X1 _13640_ (.D(net283),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[12][6] ));
 DLH_X1 _13641_ (.D(net275),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[12][7] ));
 DLH_X1 _13642_ (.D(net320),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[17][0] ));
 DLH_X1 _13643_ (.D(net310),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[17][1] ));
 DLH_X1 _13644_ (.D(net308),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[17][2] ));
 DLH_X1 _13645_ (.D(net300),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[17][3] ));
 DLH_X1 _13646_ (.D(net293),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[17][4] ));
 DLH_X1 _13647_ (.D(net287),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[17][5] ));
 DLH_X1 _13648_ (.D(net283),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[17][6] ));
 DLH_X1 _13649_ (.D(net275),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[17][7] ));
 DLH_X1 _13650_ (.D(net320),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[28][0] ));
 DLH_X1 _13651_ (.D(net310),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[28][1] ));
 DLH_X1 _13652_ (.D(net305),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[28][2] ));
 DLH_X1 _13653_ (.D(net300),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[28][3] ));
 DLH_X1 _13654_ (.D(net293),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[28][4] ));
 DLH_X1 _13655_ (.D(net287),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[28][5] ));
 DLH_X1 _13656_ (.D(net285),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[28][6] ));
 DLH_X1 _13657_ (.D(net275),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[28][7] ));
 DLH_X1 _13658_ (.D(net320),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[8][0] ));
 DLH_X1 _13659_ (.D(net310),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[8][1] ));
 DLH_X1 _13660_ (.D(net305),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[8][2] ));
 DLH_X1 _13661_ (.D(net299),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[8][3] ));
 DLH_X1 _13662_ (.D(net293),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[8][4] ));
 DLH_X1 _13663_ (.D(net287),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[8][5] ));
 DLH_X1 _13664_ (.D(net283),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[8][6] ));
 DLH_X1 _13665_ (.D(net275),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[8][7] ));
 DLH_X1 _13666_ (.D(net320),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[21][0] ));
 DLH_X1 _13667_ (.D(net310),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[21][1] ));
 DLH_X1 _13668_ (.D(net308),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[21][2] ));
 DLH_X1 _13669_ (.D(net300),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[21][3] ));
 DLH_X1 _13670_ (.D(net293),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[21][4] ));
 DLH_X1 _13671_ (.D(net287),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[21][5] ));
 DLH_X1 _13672_ (.D(net285),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[21][6] ));
 DLH_X1 _13673_ (.D(net275),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[21][7] ));
 DLH_X1 _13674_ (.D(net320),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[27][0] ));
 DLH_X1 _13675_ (.D(net310),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[27][1] ));
 DLH_X1 _13676_ (.D(net308),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[27][2] ));
 DLH_X1 _13677_ (.D(net300),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[27][3] ));
 DLH_X1 _13678_ (.D(net293),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[27][4] ));
 DLH_X1 _13679_ (.D(net287),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[27][5] ));
 DLH_X1 _13680_ (.D(net285),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[27][6] ));
 DLH_X1 _13681_ (.D(net275),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[27][7] ));
 DLH_X1 _13682_ (.D(net320),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[18][0] ));
 DLH_X1 _13683_ (.D(net310),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[18][1] ));
 DLH_X1 _13684_ (.D(net308),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[18][2] ));
 DLH_X1 _13685_ (.D(net299),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[18][3] ));
 DLH_X1 _13686_ (.D(net293),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[18][4] ));
 DLH_X1 _13687_ (.D(net287),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[18][5] ));
 DLH_X1 _13688_ (.D(net283),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[18][6] ));
 DLH_X1 _13689_ (.D(net275),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.mem[18][7] ));
 DLL_X1 _13690_ (.D(\lut.gen_sub_units_scm.__2.sub_unit_i.cg_we_global.en_i ),
    .GN(clknet_level_5_1_3218__00532_),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.cg_we_global.clk_en ));
 DLL_X1 _13691_ (.D(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__0.cg_i.en_i ),
    .GN(clknet_level_2_1_3299__00573_),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_en ));
 DLL_X1 _13692_ (.D(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__1.cg_i.en_i ),
    .GN(clknet_level_2_1_5305__00573_),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_en ));
 DLL_X1 _13693_ (.D(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__2.cg_i.en_i ),
    .GN(clknet_level_2_1_5305__00573_),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_en ));
 DLL_X1 _13694_ (.D(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__3.cg_i.en_i ),
    .GN(clknet_level_2_1_1293__00573_),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_en ));
 DLL_X1 _13695_ (.D(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__4.cg_i.en_i ),
    .GN(clknet_level_2_1_8314__00573_),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_en ));
 DLL_X1 _13696_ (.D(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__5.cg_i.en_i ),
    .GN(clknet_level_2_1_7311__00573_),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_en ));
 DLL_X1 _13697_ (.D(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__6.cg_i.en_i ),
    .GN(clknet_level_2_1_8314__00573_),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_en ));
 DLL_X1 _13698_ (.D(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__7.cg_i.en_i ),
    .GN(clknet_level_2_1_2296__00573_),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_en ));
 DLL_X1 _13699_ (.D(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__8.cg_i.en_i ),
    .GN(clknet_level_2_1_1293__00573_),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_en ));
 DLL_X1 _13700_ (.D(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__9.cg_i.en_i ),
    .GN(clknet_level_2_1_8314__00573_),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_en ));
 DLL_X1 _13701_ (.D(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__10.cg_i.en_i ),
    .GN(clknet_level_2_1_7311__00573_),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_en ));
 DLL_X1 _13702_ (.D(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__11.cg_i.en_i ),
    .GN(clknet_level_2_1_8314__00573_),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_en ));
 DLL_X1 _13703_ (.D(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__12.cg_i.en_i ),
    .GN(clknet_level_2_1_5305__00573_),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_en ));
 DLL_X1 _13704_ (.D(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__13.cg_i.en_i ),
    .GN(clknet_level_2_1_6308__00573_),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_en ));
 DLL_X1 _13705_ (.D(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__14.cg_i.en_i ),
    .GN(clknet_level_2_1_5305__00573_),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_en ));
 DLL_X1 _13706_ (.D(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__15.cg_i.en_i ),
    .GN(clknet_level_2_1_2296__00573_),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_en ));
 DLL_X1 _13707_ (.D(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__16.cg_i.en_i ),
    .GN(clknet_level_2_1_2296__00573_),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_en ));
 DLL_X1 _13708_ (.D(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__17.cg_i.en_i ),
    .GN(clknet_level_2_1_4302__00573_),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_en ));
 DLL_X1 _13709_ (.D(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__18.cg_i.en_i ),
    .GN(clknet_level_2_1_6308__00573_),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_en ));
 DLL_X1 _13710_ (.D(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__19.cg_i.en_i ),
    .GN(clknet_level_2_1_5305__00573_),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_en ));
 DLL_X1 _13711_ (.D(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__20.cg_i.en_i ),
    .GN(clknet_level_2_1_8314__00573_),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_en ));
 DLL_X1 _13712_ (.D(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__21.cg_i.en_i ),
    .GN(clknet_level_2_1_3299__00573_),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_en ));
 DLL_X1 _13713_ (.D(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__22.cg_i.en_i ),
    .GN(clknet_level_2_1_6308__00573_),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_en ));
 DLL_X1 _13714_ (.D(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__23.cg_i.en_i ),
    .GN(clknet_level_2_1_1293__00573_),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_en ));
 DLL_X1 _13715_ (.D(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__24.cg_i.en_i ),
    .GN(clknet_level_2_1_4302__00573_),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_en ));
 DLL_X1 _13716_ (.D(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__25.cg_i.en_i ),
    .GN(clknet_level_2_1_7311__00573_),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_en ));
 DLL_X1 _13717_ (.D(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__26.cg_i.en_i ),
    .GN(clknet_level_2_1_4302__00573_),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_en ));
 DLL_X1 _13718_ (.D(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__27.cg_i.en_i ),
    .GN(clknet_level_2_1_7311__00573_),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_en ));
 DLL_X1 _13719_ (.D(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__28.cg_i.en_i ),
    .GN(clknet_level_2_1_3299__00573_),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_en ));
 DLL_X1 _13720_ (.D(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__29.cg_i.en_i ),
    .GN(clknet_level_2_1_8314__00573_),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_en ));
 DLL_X1 _13721_ (.D(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__30.cg_i.en_i ),
    .GN(clknet_level_2_1_7311__00573_),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_en ));
 DLL_X1 _13722_ (.D(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__31.cg_i.en_i ),
    .GN(clknet_level_2_1_8314__00573_),
    .Q(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_en ));
 DLH_X1 _13723_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[0] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[13][0] ));
 DLH_X1 _13724_ (.D(net315),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[13][1] ));
 DLH_X1 _13725_ (.D(net309),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[13][2] ));
 DLH_X1 _13726_ (.D(net303),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[13][3] ));
 DLH_X1 _13727_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[4] ),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[13][4] ));
 DLH_X1 _13728_ (.D(net292),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[13][5] ));
 DLH_X1 _13729_ (.D(net285),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[13][6] ));
 DLH_X1 _13730_ (.D(net279),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[13][7] ));
 DLH_X1 _13731_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[0] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[1][0] ));
 DLH_X1 _13732_ (.D(net315),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[1][1] ));
 DLH_X1 _13733_ (.D(net309),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[1][2] ));
 DLH_X1 _13734_ (.D(net301),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[1][3] ));
 DLH_X1 _13735_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[4] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[1][4] ));
 DLH_X1 _13736_ (.D(net290),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[1][5] ));
 DLH_X1 _13737_ (.D(net286),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[1][6] ));
 DLH_X1 _13738_ (.D(net279),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[1][7] ));
 DLH_X1 _13739_ (.D(net319),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[26][0] ));
 DLH_X1 _13740_ (.D(net314),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[26][1] ));
 DLH_X1 _13741_ (.D(net307),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[26][2] ));
 DLH_X1 _13742_ (.D(net301),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[26][3] ));
 DLH_X1 _13743_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[4] ),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[26][4] ));
 DLH_X1 _13744_ (.D(net292),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[26][5] ));
 DLH_X1 _13745_ (.D(net285),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[26][6] ));
 DLH_X1 _13746_ (.D(net279),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[26][7] ));
 DLH_X1 _13747_ (.D(net319),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[9][0] ));
 DLH_X1 _13748_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[1] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[9][1] ));
 DLH_X1 _13749_ (.D(net309),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[9][2] ));
 DLH_X1 _13750_ (.D(net301),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[9][3] ));
 DLH_X1 _13751_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[4] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[9][4] ));
 DLH_X1 _13752_ (.D(net290),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[9][5] ));
 DLH_X1 _13753_ (.D(net286),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[9][6] ));
 DLH_X1 _13754_ (.D(net279),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[9][7] ));
 DLH_X1 _13755_ (.D(net319),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[0][0] ));
 DLH_X1 _13756_ (.D(net311),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[0][1] ));
 DLH_X1 _13757_ (.D(net306),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[0][2] ));
 DLH_X1 _13758_ (.D(net303),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[0][3] ));
 DLH_X1 _13759_ (.D(net295),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[0][4] ));
 DLH_X1 _13760_ (.D(net292),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[0][5] ));
 DLH_X1 _13761_ (.D(net285),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[0][6] ));
 DLH_X1 _13762_ (.D(net279),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[0][7] ));
 DLH_X1 _13763_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[0] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[20][0] ));
 DLH_X1 _13764_ (.D(net315),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[20][1] ));
 DLH_X1 _13765_ (.D(net306),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[20][2] ));
 DLH_X1 _13766_ (.D(net301),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[20][3] ));
 DLH_X1 _13767_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[4] ),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[20][4] ));
 DLH_X1 _13768_ (.D(net292),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[20][5] ));
 DLH_X1 _13769_ (.D(net285),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[20][6] ));
 DLH_X1 _13770_ (.D(net280),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[20][7] ));
 DLH_X1 _13771_ (.D(net319),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[2][0] ));
 DLH_X1 _13772_ (.D(net314),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[2][1] ));
 DLH_X1 _13773_ (.D(net309),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[2][2] ));
 DLH_X1 _13774_ (.D(net303),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[2][3] ));
 DLH_X1 _13775_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[4] ),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[2][4] ));
 DLH_X1 _13776_ (.D(net292),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[2][5] ));
 DLH_X1 _13777_ (.D(net285),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[2][6] ));
 DLH_X1 _13778_ (.D(net279),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[2][7] ));
 DLH_X1 _13779_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[0] ),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[25][0] ));
 DLH_X1 _13780_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[1] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[25][1] ));
 DLH_X1 _13781_ (.D(net309),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[25][2] ));
 DLH_X1 _13782_ (.D(net301),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[25][3] ));
 DLH_X1 _13783_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[4] ),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[25][4] ));
 DLH_X1 _13784_ (.D(net290),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[25][5] ));
 DLH_X1 _13785_ (.D(net286),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[25][6] ));
 DLH_X1 _13786_ (.D(net279),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[25][7] ));
 DLH_X1 _13787_ (.D(net319),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[10][0] ));
 DLH_X1 _13788_ (.D(net314),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[10][1] ));
 DLH_X1 _13789_ (.D(net307),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[10][2] ));
 DLH_X1 _13790_ (.D(net303),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[10][3] ));
 DLH_X1 _13791_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[4] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[10][4] ));
 DLH_X1 _13792_ (.D(net290),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[10][5] ));
 DLH_X1 _13793_ (.D(net286),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[10][6] ));
 DLH_X1 _13794_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[7] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[10][7] ));
 DLH_X1 _13795_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[0] ),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[3][0] ));
 DLH_X1 _13796_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[1] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[3][1] ));
 DLH_X1 _13797_ (.D(net309),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[3][2] ));
 DLH_X1 _13798_ (.D(net303),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[3][3] ));
 DLH_X1 _13799_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[4] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[3][4] ));
 DLH_X1 _13800_ (.D(net292),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[3][5] ));
 DLH_X1 _13801_ (.D(net285),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[3][6] ));
 DLH_X1 _13802_ (.D(net279),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[3][7] ));
 DLH_X1 _13803_ (.D(net319),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[16][0] ));
 DLH_X1 _13804_ (.D(net314),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[16][1] ));
 DLH_X1 _13805_ (.D(net307),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[16][2] ));
 DLH_X1 _13806_ (.D(net303),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[16][3] ));
 DLH_X1 _13807_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[4] ),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[16][4] ));
 DLH_X1 _13808_ (.D(net290),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[16][5] ));
 DLH_X1 _13809_ (.D(net285),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[16][6] ));
 DLH_X1 _13810_ (.D(net279),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[16][7] ));
 DLH_X1 _13811_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[0] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[24][0] ));
 DLH_X1 _13812_ (.D(net314),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[24][1] ));
 DLH_X1 _13813_ (.D(net307),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[24][2] ));
 DLH_X1 _13814_ (.D(net303),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[24][3] ));
 DLH_X1 _13815_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[4] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[24][4] ));
 DLH_X1 _13816_ (.D(net292),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[24][5] ));
 DLH_X1 _13817_ (.D(net285),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[24][6] ));
 DLH_X1 _13818_ (.D(net280),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[24][7] ));
 DLH_X1 _13819_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[0] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[4][0] ));
 DLH_X1 _13820_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[1] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[4][1] ));
 DLH_X1 _13821_ (.D(net307),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[4][2] ));
 DLH_X1 _13822_ (.D(net301),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[4][3] ));
 DLH_X1 _13823_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[4] ),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[4][4] ));
 DLH_X1 _13824_ (.D(net290),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[4][5] ));
 DLH_X1 _13825_ (.D(net286),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[4][6] ));
 DLH_X1 _13826_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[7] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[4][7] ));
 DLH_X1 _13827_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[0] ),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[15][0] ));
 DLH_X1 _13828_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[1] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[15][1] ));
 DLH_X1 _13829_ (.D(net307),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[15][2] ));
 DLH_X1 _13830_ (.D(net303),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[15][3] ));
 DLH_X1 _13831_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[4] ),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[15][4] ));
 DLH_X1 _13832_ (.D(net292),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[15][5] ));
 DLH_X1 _13833_ (.D(net286),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[15][6] ));
 DLH_X1 _13834_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[7] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[15][7] ));
 DLH_X1 _13835_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[0] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[11][0] ));
 DLH_X1 _13836_ (.D(net315),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[11][1] ));
 DLH_X1 _13837_ (.D(net309),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[11][2] ));
 DLH_X1 _13838_ (.D(net301),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[11][3] ));
 DLH_X1 _13839_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[4] ),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[11][4] ));
 DLH_X1 _13840_ (.D(net290),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[11][5] ));
 DLH_X1 _13841_ (.D(net286),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[11][6] ));
 DLH_X1 _13842_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[7] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[11][7] ));
 DLH_X1 _13843_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[0] ),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[5][0] ));
 DLH_X1 _13844_ (.D(net315),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[5][1] ));
 DLH_X1 _13845_ (.D(net309),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[5][2] ));
 DLH_X1 _13846_ (.D(net303),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[5][3] ));
 DLH_X1 _13847_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[4] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[5][4] ));
 DLH_X1 _13848_ (.D(net292),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[5][5] ));
 DLH_X1 _13849_ (.D(net286),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[5][6] ));
 DLH_X1 _13850_ (.D(net280),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[5][7] ));
 DLH_X1 _13851_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[0] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[23][0] ));
 DLH_X1 _13852_ (.D(net314),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[23][1] ));
 DLH_X1 _13853_ (.D(net307),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[23][2] ));
 DLH_X1 _13854_ (.D(net301),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[23][3] ));
 DLH_X1 _13855_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[4] ),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[23][4] ));
 DLH_X1 _13856_ (.D(net290),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[23][5] ));
 DLH_X1 _13857_ (.D(net286),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[23][6] ));
 DLH_X1 _13858_ (.D(net280),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[23][7] ));
 DLH_X1 _13859_ (.D(net319),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[19][0] ));
 DLH_X1 _13860_ (.D(net314),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[19][1] ));
 DLH_X1 _13861_ (.D(net307),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[19][2] ));
 DLH_X1 _13862_ (.D(net303),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[19][3] ));
 DLH_X1 _13863_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[4] ),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[19][4] ));
 DLH_X1 _13864_ (.D(net290),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[19][5] ));
 DLH_X1 _13865_ (.D(net285),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[19][6] ));
 DLH_X1 _13866_ (.D(net279),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[19][7] ));
 DLH_X1 _13867_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[0] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[31][0] ));
 DLH_X1 _13868_ (.D(net315),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[31][1] ));
 DLH_X1 _13869_ (.D(net309),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[31][2] ));
 DLH_X1 _13870_ (.D(net301),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[31][3] ));
 DLH_X1 _13871_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[4] ),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[31][4] ));
 DLH_X1 _13872_ (.D(net292),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[31][5] ));
 DLH_X1 _13873_ (.D(net285),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[31][6] ));
 DLH_X1 _13874_ (.D(net279),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[31][7] ));
 DLH_X1 _13875_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[0] ),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[6][0] ));
 DLH_X1 _13876_ (.D(net315),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[6][1] ));
 DLH_X1 _13877_ (.D(net307),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[6][2] ));
 DLH_X1 _13878_ (.D(net303),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[6][3] ));
 DLH_X1 _13879_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[4] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[6][4] ));
 DLH_X1 _13880_ (.D(net290),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[6][5] ));
 DLH_X1 _13881_ (.D(net286),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[6][6] ));
 DLH_X1 _13882_ (.D(net279),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[6][7] ));
 DLH_X1 _13883_ (.D(net319),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[14][0] ));
 DLH_X1 _13884_ (.D(net315),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[14][1] ));
 DLH_X1 _13885_ (.D(net307),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[14][2] ));
 DLH_X1 _13886_ (.D(net303),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[14][3] ));
 DLH_X1 _13887_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[4] ),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[14][4] ));
 DLH_X1 _13888_ (.D(net292),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[14][5] ));
 DLH_X1 _13889_ (.D(net285),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[14][6] ));
 DLH_X1 _13890_ (.D(net279),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[14][7] ));
 DLH_X1 _13891_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[0] ),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[30][0] ));
 DLH_X1 _13892_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[1] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[30][1] ));
 DLH_X1 _13893_ (.D(net307),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[30][2] ));
 DLH_X1 _13894_ (.D(net303),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[30][3] ));
 DLH_X1 _13895_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[4] ),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[30][4] ));
 DLH_X1 _13896_ (.D(net292),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[30][5] ));
 DLH_X1 _13897_ (.D(net286),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[30][6] ));
 DLH_X1 _13898_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[7] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[30][7] ));
 DLH_X1 _13899_ (.D(net319),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[22][0] ));
 DLH_X1 _13900_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[1] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[22][1] ));
 DLH_X1 _13901_ (.D(net309),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[22][2] ));
 DLH_X1 _13902_ (.D(net303),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[22][3] ));
 DLH_X1 _13903_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[4] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[22][4] ));
 DLH_X1 _13904_ (.D(net290),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[22][5] ));
 DLH_X1 _13905_ (.D(net285),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[22][6] ));
 DLH_X1 _13906_ (.D(net279),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[22][7] ));
 DLH_X1 _13907_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[0] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[7][0] ));
 DLH_X1 _13908_ (.D(net315),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[7][1] ));
 DLH_X1 _13909_ (.D(net309),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[7][2] ));
 DLH_X1 _13910_ (.D(net303),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[7][3] ));
 DLH_X1 _13911_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[4] ),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[7][4] ));
 DLH_X1 _13912_ (.D(net292),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[7][5] ));
 DLH_X1 _13913_ (.D(net286),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[7][6] ));
 DLH_X1 _13914_ (.D(net280),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[7][7] ));
 DLH_X1 _13915_ (.D(net319),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[29][0] ));
 DLH_X1 _13916_ (.D(net315),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[29][1] ));
 DLH_X1 _13917_ (.D(net307),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[29][2] ));
 DLH_X1 _13918_ (.D(net303),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[29][3] ));
 DLH_X1 _13919_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[4] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[29][4] ));
 DLH_X1 _13920_ (.D(net292),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[29][5] ));
 DLH_X1 _13921_ (.D(net286),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[29][6] ));
 DLH_X1 _13922_ (.D(net280),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[29][7] ));
 DLH_X1 _13923_ (.D(net319),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[12][0] ));
 DLH_X1 _13924_ (.D(net315),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[12][1] ));
 DLH_X1 _13925_ (.D(net307),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[12][2] ));
 DLH_X1 _13926_ (.D(net301),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[12][3] ));
 DLH_X1 _13927_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[4] ),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[12][4] ));
 DLH_X1 _13928_ (.D(net290),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[12][5] ));
 DLH_X1 _13929_ (.D(net285),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[12][6] ));
 DLH_X1 _13930_ (.D(net279),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[12][7] ));
 DLH_X1 _13931_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[0] ),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[17][0] ));
 DLH_X1 _13932_ (.D(net315),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[17][1] ));
 DLH_X1 _13933_ (.D(net309),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[17][2] ));
 DLH_X1 _13934_ (.D(net303),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[17][3] ));
 DLH_X1 _13935_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[4] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[17][4] ));
 DLH_X1 _13936_ (.D(net292),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[17][5] ));
 DLH_X1 _13937_ (.D(net285),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[17][6] ));
 DLH_X1 _13938_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[7] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[17][7] ));
 DLH_X1 _13939_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[0] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[28][0] ));
 DLH_X1 _13940_ (.D(net315),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[28][1] ));
 DLH_X1 _13941_ (.D(net309),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[28][2] ));
 DLH_X1 _13942_ (.D(net303),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[28][3] ));
 DLH_X1 _13943_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[4] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[28][4] ));
 DLH_X1 _13944_ (.D(net290),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[28][5] ));
 DLH_X1 _13945_ (.D(net286),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[28][6] ));
 DLH_X1 _13946_ (.D(net279),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[28][7] ));
 DLH_X1 _13947_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[0] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[8][0] ));
 DLH_X1 _13948_ (.D(net315),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[8][1] ));
 DLH_X1 _13949_ (.D(net309),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[8][2] ));
 DLH_X1 _13950_ (.D(net301),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[8][3] ));
 DLH_X1 _13951_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[4] ),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[8][4] ));
 DLH_X1 _13952_ (.D(net292),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[8][5] ));
 DLH_X1 _13953_ (.D(net285),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[8][6] ));
 DLH_X1 _13954_ (.D(net279),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[8][7] ));
 DLH_X1 _13955_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[0] ),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[21][0] ));
 DLH_X1 _13956_ (.D(net315),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[21][1] ));
 DLH_X1 _13957_ (.D(net309),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[21][2] ));
 DLH_X1 _13958_ (.D(net301),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[21][3] ));
 DLH_X1 _13959_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[4] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[21][4] ));
 DLH_X1 _13960_ (.D(net290),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[21][5] ));
 DLH_X1 _13961_ (.D(net285),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[21][6] ));
 DLH_X1 _13962_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[7] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[21][7] ));
 DLH_X1 _13963_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[0] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[27][0] ));
 DLH_X1 _13964_ (.D(net314),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[27][1] ));
 DLH_X1 _13965_ (.D(net307),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[27][2] ));
 DLH_X1 _13966_ (.D(net301),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[27][3] ));
 DLH_X1 _13967_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[4] ),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[27][4] ));
 DLH_X1 _13968_ (.D(net292),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[27][5] ));
 DLH_X1 _13969_ (.D(net286),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[27][6] ));
 DLH_X1 _13970_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[7] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[27][7] ));
 DLH_X1 _13971_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[0] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[18][0] ));
 DLH_X1 _13972_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[1] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[18][1] ));
 DLH_X1 _13973_ (.D(net307),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[18][2] ));
 DLH_X1 _13974_ (.D(net301),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[18][3] ));
 DLH_X1 _13975_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[4] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[18][4] ));
 DLH_X1 _13976_ (.D(net290),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[18][5] ));
 DLH_X1 _13977_ (.D(net286),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[18][6] ));
 DLH_X1 _13978_ (.D(net279),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.mem[18][7] ));
 DLL_X1 _13979_ (.D(\lut.gen_sub_units_scm.__1.sub_unit_i.cg_we_global.en_i ),
    .GN(clknet_level_5_1_4320__00532_),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.cg_we_global.clk_en ));
 DLL_X1 _13980_ (.D(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__0.cg_i.en_i ),
    .GN(clknet_level_2_1_2374__00576_),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_en ));
 DLL_X1 _13981_ (.D(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__1.cg_i.en_i ),
    .GN(clknet_level_2_1_7389__00576_),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_en ));
 DLL_X1 _13982_ (.D(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__2.cg_i.en_i ),
    .GN(clknet_level_2_1_1371__00576_),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_en ));
 DLL_X1 _13983_ (.D(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__3.cg_i.en_i ),
    .GN(clknet_level_2_1_7389__00576_),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_en ));
 DLL_X1 _13984_ (.D(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__4.cg_i.en_i ),
    .GN(clknet_level_2_1_8392__00576_),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_en ));
 DLL_X1 _13985_ (.D(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__5.cg_i.en_i ),
    .GN(clknet_level_2_1_7389__00576_),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_en ));
 DLL_X1 _13986_ (.D(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__6.cg_i.en_i ),
    .GN(clknet_level_2_1_7389__00576_),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_en ));
 DLL_X1 _13987_ (.D(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__7.cg_i.en_i ),
    .GN(clknet_level_2_1_6386__00576_),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_en ));
 DLL_X1 _13988_ (.D(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__8.cg_i.en_i ),
    .GN(clknet_level_2_1_6386__00576_),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_en ));
 DLL_X1 _13989_ (.D(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__9.cg_i.en_i ),
    .GN(clknet_level_2_1_3377__00576_),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_en ));
 DLL_X1 _13990_ (.D(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__10.cg_i.en_i ),
    .GN(clknet_level_2_1_3377__00576_),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_en ));
 DLL_X1 _13991_ (.D(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__11.cg_i.en_i ),
    .GN(clknet_level_2_1_8392__00576_),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_en ));
 DLL_X1 _13992_ (.D(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__12.cg_i.en_i ),
    .GN(clknet_level_2_1_2374__00576_),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_en ));
 DLL_X1 _13993_ (.D(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__13.cg_i.en_i ),
    .GN(clknet_level_2_1_5383__00576_),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_en ));
 DLL_X1 _13994_ (.D(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__14.cg_i.en_i ),
    .GN(clknet_level_2_1_2374__00576_),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_en ));
 DLL_X1 _13995_ (.D(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__15.cg_i.en_i ),
    .GN(clknet_level_2_1_5383__00576_),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_en ));
 DLL_X1 _13996_ (.D(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__16.cg_i.en_i ),
    .GN(clknet_level_2_1_4380__00576_),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_en ));
 DLL_X1 _13997_ (.D(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__17.cg_i.en_i ),
    .GN(clknet_level_2_1_6386__00576_),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_en ));
 DLL_X1 _13998_ (.D(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__18.cg_i.en_i ),
    .GN(clknet_level_2_1_4380__00576_),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_en ));
 DLL_X1 _13999_ (.D(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__19.cg_i.en_i ),
    .GN(clknet_level_2_1_4380__00576_),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_en ));
 DLL_X1 _14000_ (.D(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__20.cg_i.en_i ),
    .GN(clknet_level_2_1_5383__00576_),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_en ));
 DLL_X1 _14001_ (.D(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__21.cg_i.en_i ),
    .GN(clknet_level_2_1_6386__00576_),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_en ));
 DLL_X1 _14002_ (.D(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__22.cg_i.en_i ),
    .GN(clknet_level_2_1_1371__00576_),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_en ));
 DLL_X1 _14003_ (.D(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__23.cg_i.en_i ),
    .GN(clknet_level_2_1_4380__00576_),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_en ));
 DLL_X1 _14004_ (.D(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__24.cg_i.en_i ),
    .GN(clknet_level_2_1_6386__00576_),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_en ));
 DLL_X1 _14005_ (.D(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__25.cg_i.en_i ),
    .GN(clknet_level_2_1_4380__00576_),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_en ));
 DLL_X1 _14006_ (.D(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__26.cg_i.en_i ),
    .GN(clknet_level_2_1_1371__00576_),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_en ));
 DLL_X1 _14007_ (.D(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__27.cg_i.en_i ),
    .GN(clknet_level_2_1_8392__00576_),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_en ));
 DLL_X1 _14008_ (.D(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__28.cg_i.en_i ),
    .GN(clknet_level_2_1_8392__00576_),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_en ));
 DLL_X1 _14009_ (.D(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__29.cg_i.en_i ),
    .GN(clknet_level_2_1_8392__00576_),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_en ));
 DLL_X1 _14010_ (.D(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__30.cg_i.en_i ),
    .GN(clknet_level_2_1_8392__00576_),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_en ));
 DLL_X1 _14011_ (.D(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__31.cg_i.en_i ),
    .GN(clknet_level_2_1_5383__00576_),
    .Q(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_en ));
 DLH_X1 _14012_ (.D(net320),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[13][0] ));
 DLH_X1 _14013_ (.D(net315),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[13][1] ));
 DLH_X1 _14014_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[2] ),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[13][2] ));
 DLH_X1 _14015_ (.D(net303),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[13][3] ));
 DLH_X1 _14016_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[4] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[13][4] ));
 DLH_X1 _14017_ (.D(net292),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[13][5] ));
 DLH_X1 _14018_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[6] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[13][6] ));
 DLH_X1 _14019_ (.D(net280),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[13][7] ));
 DLH_X1 _14020_ (.D(net321),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[1][0] ));
 DLH_X1 _14021_ (.D(net315),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[1][1] ));
 DLH_X1 _14022_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[2] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[1][2] ));
 DLH_X1 _14023_ (.D(net303),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[1][3] ));
 DLH_X1 _14024_ (.D(net297),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[1][4] ));
 DLH_X1 _14025_ (.D(net292),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[1][5] ));
 DLH_X1 _14026_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[6] ),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[1][6] ));
 DLH_X1 _14027_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[7] ),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[1][7] ));
 DLH_X1 _14028_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[0] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[26][0] ));
 DLH_X1 _14029_ (.D(net315),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[26][1] ));
 DLH_X1 _14030_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[2] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[26][2] ));
 DLH_X1 _14031_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[3] ),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[26][3] ));
 DLH_X1 _14032_ (.D(net297),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[26][4] ));
 DLH_X1 _14033_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[5] ),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[26][5] ));
 DLH_X1 _14034_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[6] ),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[26][6] ));
 DLH_X1 _14035_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[7] ),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[26][7] ));
 DLH_X1 _14036_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[0] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[9][0] ));
 DLH_X1 _14037_ (.D(net315),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[9][1] ));
 DLH_X1 _14038_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[2] ),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[9][2] ));
 DLH_X1 _14039_ (.D(net303),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[9][3] ));
 DLH_X1 _14040_ (.D(net297),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[9][4] ));
 DLH_X1 _14041_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[5] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[9][5] ));
 DLH_X1 _14042_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[6] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[9][6] ));
 DLH_X1 _14043_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[7] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[9][7] ));
 DLH_X1 _14044_ (.D(net320),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[0][0] ));
 DLH_X1 _14045_ (.D(net311),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[0][1] ));
 DLH_X1 _14046_ (.D(net306),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[0][2] ));
 DLH_X1 _14047_ (.D(net303),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[0][3] ));
 DLH_X1 _14048_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[4] ),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[0][4] ));
 DLH_X1 _14049_ (.D(net292),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[0][5] ));
 DLH_X1 _14050_ (.D(net285),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[0][6] ));
 DLH_X1 _14051_ (.D(net279),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[0][7] ));
 DLH_X1 _14052_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[0] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[20][0] ));
 DLH_X1 _14053_ (.D(net315),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[20][1] ));
 DLH_X1 _14054_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[2] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[20][2] ));
 DLH_X1 _14055_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[3] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[20][3] ));
 DLH_X1 _14056_ (.D(net297),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[20][4] ));
 DLH_X1 _14057_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[5] ),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[20][5] ));
 DLH_X1 _14058_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[6] ),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[20][6] ));
 DLH_X1 _14059_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[7] ),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[20][7] ));
 DLH_X1 _14060_ (.D(net321),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[2][0] ));
 DLH_X1 _14061_ (.D(net315),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[2][1] ));
 DLH_X1 _14062_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[2] ),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[2][2] ));
 DLH_X1 _14063_ (.D(net303),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[2][3] ));
 DLH_X1 _14064_ (.D(net297),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[2][4] ));
 DLH_X1 _14065_ (.D(net292),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[2][5] ));
 DLH_X1 _14066_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[6] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[2][6] ));
 DLH_X1 _14067_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[7] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[2][7] ));
 DLH_X1 _14068_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[0] ),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[25][0] ));
 DLH_X1 _14069_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[1] ),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[25][1] ));
 DLH_X1 _14070_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[2] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[25][2] ));
 DLH_X1 _14071_ (.D(net303),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[25][3] ));
 DLH_X1 _14072_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[4] ),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[25][4] ));
 DLH_X1 _14073_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[5] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[25][5] ));
 DLH_X1 _14074_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[6] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[25][6] ));
 DLH_X1 _14075_ (.D(net280),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[25][7] ));
 DLH_X1 _14076_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[0] ),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[10][0] ));
 DLH_X1 _14077_ (.D(net315),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[10][1] ));
 DLH_X1 _14078_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[2] ),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[10][2] ));
 DLH_X1 _14079_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[3] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[10][3] ));
 DLH_X1 _14080_ (.D(net297),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[10][4] ));
 DLH_X1 _14081_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[5] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[10][5] ));
 DLH_X1 _14082_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[6] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[10][6] ));
 DLH_X1 _14083_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[7] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[10][7] ));
 DLH_X1 _14084_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[0] ),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[3][0] ));
 DLH_X1 _14085_ (.D(net315),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[3][1] ));
 DLH_X1 _14086_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[2] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[3][2] ));
 DLH_X1 _14087_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[3] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[3][3] ));
 DLH_X1 _14088_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[4] ),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[3][4] ));
 DLH_X1 _14089_ (.D(net292),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[3][5] ));
 DLH_X1 _14090_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[6] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[3][6] ));
 DLH_X1 _14091_ (.D(net280),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[3][7] ));
 DLH_X1 _14092_ (.D(net320),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[16][0] ));
 DLH_X1 _14093_ (.D(net315),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[16][1] ));
 DLH_X1 _14094_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[2] ),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[16][2] ));
 DLH_X1 _14095_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[3] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[16][3] ));
 DLH_X1 _14096_ (.D(net297),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[16][4] ));
 DLH_X1 _14097_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[5] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[16][5] ));
 DLH_X1 _14098_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[6] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[16][6] ));
 DLH_X1 _14099_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[7] ),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[16][7] ));
 DLH_X1 _14100_ (.D(net321),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[24][0] ));
 DLH_X1 _14101_ (.D(net315),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[24][1] ));
 DLH_X1 _14102_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[2] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[24][2] ));
 DLH_X1 _14103_ (.D(net303),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[24][3] ));
 DLH_X1 _14104_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[4] ),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[24][4] ));
 DLH_X1 _14105_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[5] ),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[24][5] ));
 DLH_X1 _14106_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[6] ),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[24][6] ));
 DLH_X1 _14107_ (.D(net280),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[24][7] ));
 DLH_X1 _14108_ (.D(net321),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[4][0] ));
 DLH_X1 _14109_ (.D(net315),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[4][1] ));
 DLH_X1 _14110_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[2] ),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[4][2] ));
 DLH_X1 _14111_ (.D(net303),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[4][3] ));
 DLH_X1 _14112_ (.D(net297),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[4][4] ));
 DLH_X1 _14113_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[5] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[4][5] ));
 DLH_X1 _14114_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[6] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[4][6] ));
 DLH_X1 _14115_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[7] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[4][7] ));
 DLH_X1 _14116_ (.D(net321),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[15][0] ));
 DLH_X1 _14117_ (.D(net315),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[15][1] ));
 DLH_X1 _14118_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[2] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[15][2] ));
 DLH_X1 _14119_ (.D(net303),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[15][3] ));
 DLH_X1 _14120_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[4] ),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[15][4] ));
 DLH_X1 _14121_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[5] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[15][5] ));
 DLH_X1 _14122_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[6] ),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[15][6] ));
 DLH_X1 _14123_ (.D(net280),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[15][7] ));
 DLH_X1 _14124_ (.D(net321),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[11][0] ));
 DLH_X1 _14125_ (.D(net315),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[11][1] ));
 DLH_X1 _14126_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[2] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[11][2] ));
 DLH_X1 _14127_ (.D(net303),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[11][3] ));
 DLH_X1 _14128_ (.D(net297),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[11][4] ));
 DLH_X1 _14129_ (.D(net292),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[11][5] ));
 DLH_X1 _14130_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[6] ),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[11][6] ));
 DLH_X1 _14131_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[7] ),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[11][7] ));
 DLH_X1 _14132_ (.D(net321),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[5][0] ));
 DLH_X1 _14133_ (.D(net315),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[5][1] ));
 DLH_X1 _14134_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[2] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[5][2] ));
 DLH_X1 _14135_ (.D(net303),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[5][3] ));
 DLH_X1 _14136_ (.D(net297),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[5][4] ));
 DLH_X1 _14137_ (.D(net292),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[5][5] ));
 DLH_X1 _14138_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[6] ),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[5][6] ));
 DLH_X1 _14139_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[7] ),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[5][7] ));
 DLH_X1 _14140_ (.D(net320),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[23][0] ));
 DLH_X1 _14141_ (.D(net315),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[23][1] ));
 DLH_X1 _14142_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[2] ),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[23][2] ));
 DLH_X1 _14143_ (.D(net303),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[23][3] ));
 DLH_X1 _14144_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[4] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[23][4] ));
 DLH_X1 _14145_ (.D(net292),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[23][5] ));
 DLH_X1 _14146_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[6] ),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[23][6] ));
 DLH_X1 _14147_ (.D(net280),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[23][7] ));
 DLH_X1 _14148_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[0] ),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[19][0] ));
 DLH_X1 _14149_ (.D(net315),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[19][1] ));
 DLH_X1 _14150_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[2] ),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[19][2] ));
 DLH_X1 _14151_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[3] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[19][3] ));
 DLH_X1 _14152_ (.D(net297),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[19][4] ));
 DLH_X1 _14153_ (.D(net292),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[19][5] ));
 DLH_X1 _14154_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[6] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[19][6] ));
 DLH_X1 _14155_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[7] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[19][7] ));
 DLH_X1 _14156_ (.D(net321),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[31][0] ));
 DLH_X1 _14157_ (.D(net315),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[31][1] ));
 DLH_X1 _14158_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[2] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[31][2] ));
 DLH_X1 _14159_ (.D(net303),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[31][3] ));
 DLH_X1 _14160_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[4] ),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[31][4] ));
 DLH_X1 _14161_ (.D(net292),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[31][5] ));
 DLH_X1 _14162_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[6] ),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[31][6] ));
 DLH_X1 _14163_ (.D(net280),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[31][7] ));
 DLH_X1 _14164_ (.D(net321),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[6][0] ));
 DLH_X1 _14165_ (.D(net315),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[6][1] ));
 DLH_X1 _14166_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[2] ),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[6][2] ));
 DLH_X1 _14167_ (.D(net303),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[6][3] ));
 DLH_X1 _14168_ (.D(net297),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[6][4] ));
 DLH_X1 _14169_ (.D(net292),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[6][5] ));
 DLH_X1 _14170_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[6] ),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[6][6] ));
 DLH_X1 _14171_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[7] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[6][7] ));
 DLH_X1 _14172_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[0] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[14][0] ));
 DLH_X1 _14173_ (.D(net315),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[14][1] ));
 DLH_X1 _14174_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[2] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[14][2] ));
 DLH_X1 _14175_ (.D(net303),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[14][3] ));
 DLH_X1 _14176_ (.D(net297),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[14][4] ));
 DLH_X1 _14177_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[5] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[14][5] ));
 DLH_X1 _14178_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[6] ),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[14][6] ));
 DLH_X1 _14179_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[7] ),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[14][7] ));
 DLH_X1 _14180_ (.D(net320),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[30][0] ));
 DLH_X1 _14181_ (.D(net315),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[30][1] ));
 DLH_X1 _14182_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[2] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[30][2] ));
 DLH_X1 _14183_ (.D(net303),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[30][3] ));
 DLH_X1 _14184_ (.D(net297),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[30][4] ));
 DLH_X1 _14185_ (.D(net292),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[30][5] ));
 DLH_X1 _14186_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[6] ),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[30][6] ));
 DLH_X1 _14187_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[7] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[30][7] ));
 DLH_X1 _14188_ (.D(net321),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[22][0] ));
 DLH_X1 _14189_ (.D(net315),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[22][1] ));
 DLH_X1 _14190_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[2] ),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[22][2] ));
 DLH_X1 _14191_ (.D(net303),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[22][3] ));
 DLH_X1 _14192_ (.D(net297),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[22][4] ));
 DLH_X1 _14193_ (.D(net292),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[22][5] ));
 DLH_X1 _14194_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[6] ),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[22][6] ));
 DLH_X1 _14195_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[7] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[22][7] ));
 DLH_X1 _14196_ (.D(net321),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[7][0] ));
 DLH_X1 _14197_ (.D(net315),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[7][1] ));
 DLH_X1 _14198_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[2] ),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[7][2] ));
 DLH_X1 _14199_ (.D(net303),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[7][3] ));
 DLH_X1 _14200_ (.D(net297),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[7][4] ));
 DLH_X1 _14201_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[5] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[7][5] ));
 DLH_X1 _14202_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[6] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[7][6] ));
 DLH_X1 _14203_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[7] ),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[7][7] ));
 DLH_X1 _14204_ (.D(net321),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[29][0] ));
 DLH_X1 _14205_ (.D(net315),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[29][1] ));
 DLH_X1 _14206_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[2] ),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[29][2] ));
 DLH_X1 _14207_ (.D(net303),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[29][3] ));
 DLH_X1 _14208_ (.D(net297),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[29][4] ));
 DLH_X1 _14209_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[5] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[29][5] ));
 DLH_X1 _14210_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[6] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[29][6] ));
 DLH_X1 _14211_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[7] ),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[29][7] ));
 DLH_X1 _14212_ (.D(net321),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[12][0] ));
 DLH_X1 _14213_ (.D(net315),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[12][1] ));
 DLH_X1 _14214_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[2] ),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[12][2] ));
 DLH_X1 _14215_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[3] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[12][3] ));
 DLH_X1 _14216_ (.D(net297),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[12][4] ));
 DLH_X1 _14217_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[5] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[12][5] ));
 DLH_X1 _14218_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[6] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[12][6] ));
 DLH_X1 _14219_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[7] ),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[12][7] ));
 DLH_X1 _14220_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[0] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[17][0] ));
 DLH_X1 _14221_ (.D(net315),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[17][1] ));
 DLH_X1 _14222_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[2] ),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[17][2] ));
 DLH_X1 _14223_ (.D(net303),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[17][3] ));
 DLH_X1 _14224_ (.D(net297),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[17][4] ));
 DLH_X1 _14225_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[5] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[17][5] ));
 DLH_X1 _14226_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[6] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[17][6] ));
 DLH_X1 _14227_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[7] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[17][7] ));
 DLH_X1 _14228_ (.D(net321),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[28][0] ));
 DLH_X1 _14229_ (.D(net315),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[28][1] ));
 DLH_X1 _14230_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[2] ),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[28][2] ));
 DLH_X1 _14231_ (.D(net303),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[28][3] ));
 DLH_X1 _14232_ (.D(net297),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[28][4] ));
 DLH_X1 _14233_ (.D(net292),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[28][5] ));
 DLH_X1 _14234_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[6] ),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[28][6] ));
 DLH_X1 _14235_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[7] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[28][7] ));
 DLH_X1 _14236_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[0] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[8][0] ));
 DLH_X1 _14237_ (.D(net315),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[8][1] ));
 DLH_X1 _14238_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[2] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[8][2] ));
 DLH_X1 _14239_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[3] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[8][3] ));
 DLH_X1 _14240_ (.D(net297),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[8][4] ));
 DLH_X1 _14241_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[5] ),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[8][5] ));
 DLH_X1 _14242_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[6] ),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[8][6] ));
 DLH_X1 _14243_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[7] ),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[8][7] ));
 DLH_X1 _14244_ (.D(net321),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[21][0] ));
 DLH_X1 _14245_ (.D(net315),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[21][1] ));
 DLH_X1 _14246_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[2] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[21][2] ));
 DLH_X1 _14247_ (.D(net303),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[21][3] ));
 DLH_X1 _14248_ (.D(net297),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[21][4] ));
 DLH_X1 _14249_ (.D(net292),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[21][5] ));
 DLH_X1 _14250_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[6] ),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[21][6] ));
 DLH_X1 _14251_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[7] ),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[21][7] ));
 DLH_X1 _14252_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[0] ),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[27][0] ));
 DLH_X1 _14253_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[1] ),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[27][1] ));
 DLH_X1 _14254_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[2] ),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[27][2] ));
 DLH_X1 _14255_ (.D(net303),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[27][3] ));
 DLH_X1 _14256_ (.D(net297),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[27][4] ));
 DLH_X1 _14257_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[5] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[27][5] ));
 DLH_X1 _14258_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[6] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[27][6] ));
 DLH_X1 _14259_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[7] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[27][7] ));
 DLH_X1 _14260_ (.D(net321),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[18][0] ));
 DLH_X1 _14261_ (.D(net315),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[18][1] ));
 DLH_X1 _14262_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[2] ),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[18][2] ));
 DLH_X1 _14263_ (.D(net303),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[18][3] ));
 DLH_X1 _14264_ (.D(net297),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[18][4] ));
 DLH_X1 _14265_ (.D(net292),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[18][5] ));
 DLH_X1 _14266_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[6] ),
    .G(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[18][6] ));
 DLH_X1 _14267_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[7] ),
    .G(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.mem[18][7] ));
 DLL_X1 _14268_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.cg_we_global.en_i ),
    .GN(clknet_level_5_1_4320__00532_),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.cg_we_global.clk_en ));
 DLL_X1 _14269_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__0.cg_i.en_i ),
    .GN(clknet_level_2_1_5407__00579_),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_en ));
 DLL_X1 _14270_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__1.cg_i.en_i ),
    .GN(clknet_level_2_1_5407__00579_),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_en ));
 DLL_X1 _14271_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__2.cg_i.en_i ),
    .GN(clknet_level_2_1_1395__00579_),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_en ));
 DLL_X1 _14272_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__3.cg_i.en_i ),
    .GN(clknet_level_2_1_7413__00579_),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_en ));
 DLL_X1 _14273_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__4.cg_i.en_i ),
    .GN(clknet_level_2_1_5407__00579_),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_en ));
 DLL_X1 _14274_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__5.cg_i.en_i ),
    .GN(clknet_level_2_1_4404__00579_),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_en ));
 DLL_X1 _14275_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__6.cg_i.en_i ),
    .GN(clknet_level_2_1_5407__00579_),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_en ));
 DLL_X1 _14276_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__7.cg_i.en_i ),
    .GN(clknet_level_2_1_8416__00579_),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_en ));
 DLL_X1 _14277_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__8.cg_i.en_i ),
    .GN(clknet_level_2_1_7413__00579_),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_en ));
 DLL_X1 _14278_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__9.cg_i.en_i ),
    .GN(clknet_level_2_1_3401__00579_),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_en ));
 DLL_X1 _14279_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__10.cg_i.en_i ),
    .GN(clknet_level_2_1_7413__00579_),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_en ));
 DLL_X1 _14280_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__11.cg_i.en_i ),
    .GN(clknet_level_2_1_8416__00579_),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_en ));
 DLL_X1 _14281_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__12.cg_i.en_i ),
    .GN(clknet_level_2_1_1395__00579_),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_en ));
 DLL_X1 _14282_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__13.cg_i.en_i ),
    .GN(clknet_level_2_1_6410__00579_),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_en ));
 DLL_X1 _14283_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__14.cg_i.en_i ),
    .GN(clknet_level_2_1_3401__00579_),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_en ));
 DLL_X1 _14284_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__15.cg_i.en_i ),
    .GN(clknet_level_2_1_8416__00579_),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_en ));
 DLL_X1 _14285_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__16.cg_i.en_i ),
    .GN(clknet_level_2_1_3401__00579_),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_en ));
 DLL_X1 _14286_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__17.cg_i.en_i ),
    .GN(clknet_level_2_1_8416__00579_),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_en ));
 DLL_X1 _14287_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__18.cg_i.en_i ),
    .GN(clknet_level_2_1_6410__00579_),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_en ));
 DLL_X1 _14288_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__19.cg_i.en_i ),
    .GN(clknet_level_2_1_4404__00579_),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_en ));
 DLL_X1 _14289_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__20.cg_i.en_i ),
    .GN(clknet_level_2_1_8416__00579_),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_en ));
 DLL_X1 _14290_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__21.cg_i.en_i ),
    .GN(clknet_level_2_1_4404__00579_),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_en ));
 DLL_X1 _14291_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__22.cg_i.en_i ),
    .GN(clknet_level_2_1_2398__00579_),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_en ));
 DLL_X1 _14292_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__23.cg_i.en_i ),
    .GN(clknet_level_2_1_6410__00579_),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_en ));
 DLL_X1 _14293_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__24.cg_i.en_i ),
    .GN(clknet_level_2_1_1395__00579_),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_en ));
 DLL_X1 _14294_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__25.cg_i.en_i ),
    .GN(clknet_level_2_1_6410__00579_),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_en ));
 DLL_X1 _14295_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__26.cg_i.en_i ),
    .GN(clknet_level_2_1_7413__00579_),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_en ));
 DLL_X1 _14296_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__27.cg_i.en_i ),
    .GN(clknet_level_2_1_7413__00579_),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_en ));
 DLL_X1 _14297_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__28.cg_i.en_i ),
    .GN(clknet_level_2_1_4404__00579_),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_en ));
 DLL_X1 _14298_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__29.cg_i.en_i ),
    .GN(clknet_level_2_1_4404__00579_),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_en ));
 DLL_X1 _14299_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__30.cg_i.en_i ),
    .GN(clknet_level_2_1_4404__00579_),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_en ));
 DLL_X1 _14300_ (.D(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__31.cg_i.en_i ),
    .GN(clknet_level_2_1_6410__00579_),
    .Q(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_en ));
 DLL_X1 _14301_ (.D(net29),
    .GN(clknet_level_8_1_18_clk_i),
    .Q(\lut.cg_we_global.clk_en ));
 BUF_X4 wire232 (.A(net237),
    .Z(net232));
 BUF_X4 max_cap233 (.A(net236),
    .Z(net233));
 BUF_X4 wire234 (.A(net235),
    .Z(net234));
 BUF_X8 max_cap235 (.A(net236),
    .Z(net235));
 BUF_X4 wire236 (.A(net237),
    .Z(net236));
 BUF_X8 max_cap237 (.A(_00993_),
    .Z(net237));
 BUF_X8 max_cap238 (.A(net239),
    .Z(net238));
 BUF_X8 max_cap239 (.A(_00989_),
    .Z(net239));
 BUF_X8 max_cap240 (.A(net242),
    .Z(net240));
 BUF_X16 max_cap241 (.A(net242),
    .Z(net241));
 BUF_X16 max_cap242 (.A(net243),
    .Z(net242));
 BUF_X8 wire243 (.A(_00989_),
    .Z(net243));
 BUF_X4 max_cap244 (.A(_00986_),
    .Z(net244));
 BUF_X4 max_cap245 (.A(_00986_),
    .Z(net245));
 BUF_X4 wire246 (.A(_00986_),
    .Z(net246));
 BUF_X4 max_cap247 (.A(net249),
    .Z(net247));
 BUF_X8 max_cap248 (.A(net252),
    .Z(net248));
 BUF_X8 max_cap249 (.A(net252),
    .Z(net249));
 BUF_X4 wire250 (.A(net251),
    .Z(net250));
 BUF_X8 max_cap251 (.A(net252),
    .Z(net251));
 BUF_X8 max_cap252 (.A(_00986_),
    .Z(net252));
 BUF_X4 max_cap253 (.A(_00975_),
    .Z(net253));
 BUF_X8 max_cap254 (.A(net255),
    .Z(net254));
 BUF_X4 max_cap255 (.A(net260),
    .Z(net255));
 BUF_X4 max_cap256 (.A(net260),
    .Z(net256));
 BUF_X4 max_cap257 (.A(net259),
    .Z(net257));
 BUF_X8 max_cap258 (.A(net259),
    .Z(net258));
 BUF_X8 max_cap259 (.A(net260),
    .Z(net259));
 BUF_X4 wire260 (.A(_00975_),
    .Z(net260));
 BUF_X4 max_cap261 (.A(net262),
    .Z(net261));
 BUF_X4 max_cap262 (.A(_00975_),
    .Z(net262));
 BUF_X16 max_cap263 (.A(net265),
    .Z(net263));
 BUF_X16 max_length264 (.A(net265),
    .Z(net264));
 BUF_X16 max_cap265 (.A(_00964_),
    .Z(net265));
 BUF_X8 max_cap266 (.A(net272),
    .Z(net266));
 BUF_X4 max_cap267 (.A(net268),
    .Z(net267));
 BUF_X4 max_cap268 (.A(net269),
    .Z(net268));
 BUF_X4 wire269 (.A(net271),
    .Z(net269));
 BUF_X4 max_cap270 (.A(net271),
    .Z(net270));
 BUF_X4 max_cap271 (.A(_00950_),
    .Z(net271));
 BUF_X4 max_cap272 (.A(_00950_),
    .Z(net272));
 BUF_X4 wire273 (.A(net274),
    .Z(net273));
 BUF_X4 wire274 (.A(_00950_),
    .Z(net274));
 BUF_X16 wire275 (.A(net277),
    .Z(net275));
 BUF_X16 max_cap276 (.A(net277),
    .Z(net276));
 BUF_X16 max_cap277 (.A(net280),
    .Z(net277));
 BUF_X16 max_cap278 (.A(net279),
    .Z(net278));
 BUF_X16 max_cap279 (.A(net280),
    .Z(net279));
 BUF_X16 max_cap280 (.A(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[7] ),
    .Z(net280));
 BUF_X16 max_cap281 (.A(net286),
    .Z(net281));
 BUF_X16 max_cap282 (.A(net284),
    .Z(net282));
 BUF_X16 max_cap283 (.A(net285),
    .Z(net283));
 BUF_X16 max_cap284 (.A(net285),
    .Z(net284));
 BUF_X16 max_cap285 (.A(net286),
    .Z(net285));
 BUF_X16 max_cap286 (.A(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[6] ),
    .Z(net286));
 BUF_X32 max_cap287 (.A(net288),
    .Z(net287));
 BUF_X16 wire288 (.A(net292),
    .Z(net288));
 BUF_X16 max_cap289 (.A(net290),
    .Z(net289));
 BUF_X16 max_cap290 (.A(net292),
    .Z(net290));
 BUF_X16 max_cap291 (.A(net292),
    .Z(net291));
 BUF_X16 wire292 (.A(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[5] ),
    .Z(net292));
 BUF_X16 max_cap293 (.A(net297),
    .Z(net293));
 BUF_X32 max_cap294 (.A(net295),
    .Z(net294));
 BUF_X16 wire295 (.A(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[4] ),
    .Z(net295));
 BUF_X16 max_cap296 (.A(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[4] ),
    .Z(net296));
 BUF_X16 max_cap297 (.A(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[4] ),
    .Z(net297));
 BUF_X16 max_cap298 (.A(net303),
    .Z(net298));
 BUF_X16 max_cap299 (.A(net300),
    .Z(net299));
 BUF_X16 max_cap300 (.A(net303),
    .Z(net300));
 BUF_X16 max_cap301 (.A(net303),
    .Z(net301));
 BUF_X16 max_cap302 (.A(net303),
    .Z(net302));
 BUF_X16 max_cap303 (.A(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[3] ),
    .Z(net303));
 BUF_X16 max_cap304 (.A(net307),
    .Z(net304));
 BUF_X16 max_cap305 (.A(net306),
    .Z(net305));
 BUF_X16 max_cap306 (.A(net307),
    .Z(net306));
 BUF_X16 max_cap307 (.A(net309),
    .Z(net307));
 BUF_X16 max_cap308 (.A(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[2] ),
    .Z(net308));
 BUF_X16 max_cap309 (.A(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[2] ),
    .Z(net309));
 BUF_X16 wire310 (.A(net315),
    .Z(net310));
 BUF_X16 max_cap311 (.A(net315),
    .Z(net311));
 BUF_X16 max_cap312 (.A(net313),
    .Z(net312));
 BUF_X16 max_cap313 (.A(net314),
    .Z(net313));
 BUF_X16 wire314 (.A(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[1] ),
    .Z(net314));
 BUF_X16 max_cap315 (.A(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[1] ),
    .Z(net315));
 BUF_X16 max_cap316 (.A(net317),
    .Z(net316));
 BUF_X16 max_cap317 (.A(net319),
    .Z(net317));
 BUF_X16 max_cap318 (.A(net319),
    .Z(net318));
 BUF_X16 wire319 (.A(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[0] ),
    .Z(net319));
 BUF_X16 max_cap320 (.A(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[0] ),
    .Z(net320));
 BUF_X16 max_cap321 (.A(\lut.gen_sub_units_scm.__0.sub_unit_i.wdata_a_i[0] ),
    .Z(net321));
 BUF_X4 clkbuf_0_clk_i (.A(clk_i),
    .Z(clknet_0_clk_i));
 BUF_X4 clkbuf_3_0__f_clk_i (.A(clknet_0_clk_i),
    .Z(clknet_3_0__leaf_clk_i));
 BUF_X4 clkbuf_3_1__f_clk_i (.A(clknet_0_clk_i),
    .Z(clknet_3_1__leaf_clk_i));
 BUF_X4 clkbuf_3_2__f_clk_i (.A(clknet_0_clk_i),
    .Z(clknet_3_2__leaf_clk_i));
 BUF_X4 clkbuf_3_3__f_clk_i (.A(clknet_0_clk_i),
    .Z(clknet_3_3__leaf_clk_i));
 BUF_X4 clkbuf_3_4__f_clk_i (.A(clknet_0_clk_i),
    .Z(clknet_3_4__leaf_clk_i));
 BUF_X4 clkbuf_3_5__f_clk_i (.A(clknet_0_clk_i),
    .Z(clknet_3_5__leaf_clk_i));
 BUF_X4 clkbuf_3_6__f_clk_i (.A(clknet_0_clk_i),
    .Z(clknet_3_6__leaf_clk_i));
 BUF_X4 clkbuf_3_7__f_clk_i (.A(clknet_0_clk_i),
    .Z(clknet_3_7__leaf_clk_i));
 BUF_X4 clkbuf_level_0_1_10_clk_i (.A(clknet_3_0__leaf_clk_i),
    .Z(clknet_level_0_1_10_clk_i));
 BUF_X4 clkbuf_level_1_1_11_clk_i (.A(clknet_level_0_1_10_clk_i),
    .Z(clknet_level_1_1_11_clk_i));
 BUF_X4 clkbuf_level_2_1_12_clk_i (.A(clknet_level_1_1_11_clk_i),
    .Z(clknet_level_2_1_12_clk_i));
 BUF_X4 clkbuf_level_3_1_13_clk_i (.A(clknet_level_2_1_12_clk_i),
    .Z(clknet_level_3_1_13_clk_i));
 BUF_X4 clkbuf_level_4_1_14_clk_i (.A(clknet_level_3_1_13_clk_i),
    .Z(clknet_level_4_1_14_clk_i));
 BUF_X4 clkbuf_level_5_1_15_clk_i (.A(clknet_level_4_1_14_clk_i),
    .Z(clknet_level_5_1_15_clk_i));
 BUF_X4 clkbuf_level_6_1_16_clk_i (.A(clknet_level_5_1_15_clk_i),
    .Z(clknet_level_6_1_16_clk_i));
 BUF_X4 clkbuf_level_7_1_17_clk_i (.A(clknet_level_6_1_16_clk_i),
    .Z(clknet_level_7_1_17_clk_i));
 BUF_X4 clkbuf_level_8_1_18_clk_i (.A(clknet_level_7_1_17_clk_i),
    .Z(clknet_level_8_1_18_clk_i));
 BUF_X4 clkbuf_level_0_1_2417_clk_i (.A(clknet_3_1__leaf_clk_i),
    .Z(clknet_level_0_1_2417_clk_i));
 BUF_X4 clkbuf_level_1_1_2418_clk_i (.A(clknet_level_0_1_2417_clk_i),
    .Z(clknet_level_1_1_2418_clk_i));
 BUF_X4 clkbuf_level_2_1_2419_clk_i (.A(clknet_level_1_1_2418_clk_i),
    .Z(clknet_level_2_1_2419_clk_i));
 BUF_X4 clkbuf_level_3_1_2420_clk_i (.A(clknet_level_2_1_2419_clk_i),
    .Z(clknet_level_3_1_2420_clk_i));
 BUF_X4 clkbuf_level_4_1_2421_clk_i (.A(clknet_level_3_1_2420_clk_i),
    .Z(clknet_level_4_1_2421_clk_i));
 BUF_X4 clkbuf_level_5_1_2422_clk_i (.A(clknet_level_4_1_2421_clk_i),
    .Z(clknet_level_5_1_2422_clk_i));
 BUF_X4 clkbuf_level_6_1_2423_clk_i (.A(clknet_level_5_1_2422_clk_i),
    .Z(clknet_level_6_1_2423_clk_i));
 BUF_X4 clkbuf_level_7_1_2424_clk_i (.A(clknet_level_6_1_2423_clk_i),
    .Z(clknet_level_7_1_2424_clk_i));
 BUF_X4 clkbuf_level_8_1_2425_clk_i (.A(clknet_level_7_1_2424_clk_i),
    .Z(clknet_level_8_1_2425_clk_i));
 BUF_X4 clkbuf_level_0_1_3426_clk_i (.A(clknet_3_2__leaf_clk_i),
    .Z(clknet_level_0_1_3426_clk_i));
 BUF_X4 clkbuf_level_1_1_3427_clk_i (.A(clknet_level_0_1_3426_clk_i),
    .Z(clknet_level_1_1_3427_clk_i));
 BUF_X4 clkbuf_level_2_1_3428_clk_i (.A(clknet_level_1_1_3427_clk_i),
    .Z(clknet_level_2_1_3428_clk_i));
 BUF_X4 clkbuf_level_3_1_3429_clk_i (.A(clknet_level_2_1_3428_clk_i),
    .Z(clknet_level_3_1_3429_clk_i));
 BUF_X4 clkbuf_level_4_1_3430_clk_i (.A(clknet_level_3_1_3429_clk_i),
    .Z(clknet_level_4_1_3430_clk_i));
 BUF_X4 clkbuf_level_5_1_3431_clk_i (.A(clknet_level_4_1_3430_clk_i),
    .Z(clknet_level_5_1_3431_clk_i));
 BUF_X4 clkbuf_level_6_1_3432_clk_i (.A(clknet_level_5_1_3431_clk_i),
    .Z(clknet_level_6_1_3432_clk_i));
 BUF_X4 clkbuf_level_7_1_3433_clk_i (.A(clknet_level_6_1_3432_clk_i),
    .Z(clknet_level_7_1_3433_clk_i));
 BUF_X4 clkbuf_level_8_1_3434_clk_i (.A(clknet_level_7_1_3433_clk_i),
    .Z(clknet_level_8_1_3434_clk_i));
 BUF_X4 clkbuf_level_0_1_4435_clk_i (.A(clknet_3_3__leaf_clk_i),
    .Z(clknet_level_0_1_4435_clk_i));
 BUF_X4 clkbuf_level_1_1_4436_clk_i (.A(clknet_level_0_1_4435_clk_i),
    .Z(clknet_level_1_1_4436_clk_i));
 BUF_X4 clkbuf_level_2_1_4437_clk_i (.A(clknet_level_1_1_4436_clk_i),
    .Z(clknet_level_2_1_4437_clk_i));
 BUF_X4 clkbuf_level_3_1_4438_clk_i (.A(clknet_level_2_1_4437_clk_i),
    .Z(clknet_level_3_1_4438_clk_i));
 BUF_X4 clkbuf_level_4_1_4439_clk_i (.A(clknet_level_3_1_4438_clk_i),
    .Z(clknet_level_4_1_4439_clk_i));
 BUF_X4 clkbuf_level_5_1_4440_clk_i (.A(clknet_level_4_1_4439_clk_i),
    .Z(clknet_level_5_1_4440_clk_i));
 BUF_X4 clkbuf_level_6_1_4441_clk_i (.A(clknet_level_5_1_4440_clk_i),
    .Z(clknet_level_6_1_4441_clk_i));
 BUF_X4 clkbuf_level_7_1_4442_clk_i (.A(clknet_level_6_1_4441_clk_i),
    .Z(clknet_level_7_1_4442_clk_i));
 BUF_X4 clkbuf_level_8_1_4443_clk_i (.A(clknet_level_7_1_4442_clk_i),
    .Z(clknet_level_8_1_4443_clk_i));
 BUF_X4 clkbuf_level_0_1_5444_clk_i (.A(clknet_3_4__leaf_clk_i),
    .Z(clknet_level_0_1_5444_clk_i));
 BUF_X4 clkbuf_level_1_1_5445_clk_i (.A(clknet_level_0_1_5444_clk_i),
    .Z(clknet_level_1_1_5445_clk_i));
 BUF_X4 clkbuf_level_2_1_5446_clk_i (.A(clknet_level_1_1_5445_clk_i),
    .Z(clknet_level_2_1_5446_clk_i));
 BUF_X4 clkbuf_level_3_1_5447_clk_i (.A(clknet_level_2_1_5446_clk_i),
    .Z(clknet_level_3_1_5447_clk_i));
 BUF_X4 clkbuf_level_4_1_5448_clk_i (.A(clknet_level_3_1_5447_clk_i),
    .Z(clknet_level_4_1_5448_clk_i));
 BUF_X4 clkbuf_level_5_1_5449_clk_i (.A(clknet_level_4_1_5448_clk_i),
    .Z(clknet_level_5_1_5449_clk_i));
 BUF_X4 clkbuf_level_6_1_5450_clk_i (.A(clknet_level_5_1_5449_clk_i),
    .Z(clknet_level_6_1_5450_clk_i));
 BUF_X4 clkbuf_level_7_1_5451_clk_i (.A(clknet_level_6_1_5450_clk_i),
    .Z(clknet_level_7_1_5451_clk_i));
 BUF_X4 clkbuf_level_8_1_5452_clk_i (.A(clknet_level_7_1_5451_clk_i),
    .Z(clknet_level_8_1_5452_clk_i));
 BUF_X4 clkbuf_level_0_1_6453_clk_i (.A(clknet_3_5__leaf_clk_i),
    .Z(clknet_level_0_1_6453_clk_i));
 BUF_X4 clkbuf_level_1_1_6454_clk_i (.A(clknet_level_0_1_6453_clk_i),
    .Z(clknet_level_1_1_6454_clk_i));
 BUF_X4 clkbuf_level_2_1_6455_clk_i (.A(clknet_level_1_1_6454_clk_i),
    .Z(clknet_level_2_1_6455_clk_i));
 BUF_X4 clkbuf_level_3_1_6456_clk_i (.A(clknet_level_2_1_6455_clk_i),
    .Z(clknet_level_3_1_6456_clk_i));
 BUF_X4 clkbuf_level_4_1_6457_clk_i (.A(clknet_level_3_1_6456_clk_i),
    .Z(clknet_level_4_1_6457_clk_i));
 BUF_X4 clkbuf_level_5_1_6458_clk_i (.A(clknet_level_4_1_6457_clk_i),
    .Z(clknet_level_5_1_6458_clk_i));
 BUF_X4 clkbuf_level_6_1_6459_clk_i (.A(clknet_level_5_1_6458_clk_i),
    .Z(clknet_level_6_1_6459_clk_i));
 BUF_X4 clkbuf_level_7_1_6460_clk_i (.A(clknet_level_6_1_6459_clk_i),
    .Z(clknet_level_7_1_6460_clk_i));
 BUF_X4 clkbuf_level_8_1_6461_clk_i (.A(clknet_level_7_1_6460_clk_i),
    .Z(clknet_level_8_1_6461_clk_i));
 BUF_X4 clkbuf_level_0_1_7462_clk_i (.A(clknet_3_6__leaf_clk_i),
    .Z(clknet_level_0_1_7462_clk_i));
 BUF_X4 clkbuf_level_1_1_7463_clk_i (.A(clknet_level_0_1_7462_clk_i),
    .Z(clknet_level_1_1_7463_clk_i));
 BUF_X4 clkbuf_level_2_1_7464_clk_i (.A(clknet_level_1_1_7463_clk_i),
    .Z(clknet_level_2_1_7464_clk_i));
 BUF_X4 clkbuf_level_3_1_7465_clk_i (.A(clknet_level_2_1_7464_clk_i),
    .Z(clknet_level_3_1_7465_clk_i));
 BUF_X4 clkbuf_level_4_1_7466_clk_i (.A(clknet_level_3_1_7465_clk_i),
    .Z(clknet_level_4_1_7466_clk_i));
 BUF_X4 clkbuf_level_5_1_7467_clk_i (.A(clknet_level_4_1_7466_clk_i),
    .Z(clknet_level_5_1_7467_clk_i));
 BUF_X4 clkbuf_level_6_1_7468_clk_i (.A(clknet_level_5_1_7467_clk_i),
    .Z(clknet_level_6_1_7468_clk_i));
 BUF_X4 clkbuf_level_7_1_7469_clk_i (.A(clknet_level_6_1_7468_clk_i),
    .Z(clknet_level_7_1_7469_clk_i));
 BUF_X4 clkbuf_level_8_1_7470_clk_i (.A(clknet_level_7_1_7469_clk_i),
    .Z(clknet_level_8_1_7470_clk_i));
 BUF_X4 clkbuf_level_0_1_8471_clk_i (.A(clknet_3_7__leaf_clk_i),
    .Z(clknet_level_0_1_8471_clk_i));
 BUF_X4 clkbuf_level_1_1_8472_clk_i (.A(clknet_level_0_1_8471_clk_i),
    .Z(clknet_level_1_1_8472_clk_i));
 BUF_X4 clkbuf_level_2_1_8473_clk_i (.A(clknet_level_1_1_8472_clk_i),
    .Z(clknet_level_2_1_8473_clk_i));
 BUF_X4 clkbuf_level_3_1_8474_clk_i (.A(clknet_level_2_1_8473_clk_i),
    .Z(clknet_level_3_1_8474_clk_i));
 BUF_X4 clkbuf_level_4_1_8475_clk_i (.A(clknet_level_3_1_8474_clk_i),
    .Z(clknet_level_4_1_8475_clk_i));
 BUF_X4 clkbuf_level_5_1_8476_clk_i (.A(clknet_level_4_1_8475_clk_i),
    .Z(clknet_level_5_1_8476_clk_i));
 BUF_X4 clkbuf_level_6_1_8477_clk_i (.A(clknet_level_5_1_8476_clk_i),
    .Z(clknet_level_6_1_8477_clk_i));
 BUF_X4 clkbuf_level_7_1_8478_clk_i (.A(clknet_level_6_1_8477_clk_i),
    .Z(clknet_level_7_1_8478_clk_i));
 BUF_X4 clkbuf_level_8_1_8479_clk_i (.A(clknet_level_7_1_8478_clk_i),
    .Z(clknet_level_8_1_8479_clk_i));
 BUF_X4 clkbuf_0__00532_ (.A(_00532_),
    .Z(clknet_0__00532_));
 BUF_X4 clkbuf_2_0__f__00532_ (.A(clknet_0__00532_),
    .Z(clknet_2_0__leaf__00532_));
 BUF_X4 clkbuf_2_1__f__00532_ (.A(clknet_0__00532_),
    .Z(clknet_2_1__leaf__00532_));
 BUF_X4 clkbuf_2_2__f__00532_ (.A(clknet_0__00532_),
    .Z(clknet_2_2__leaf__00532_));
 BUF_X4 clkbuf_2_3__f__00532_ (.A(clknet_0__00532_),
    .Z(clknet_2_3__leaf__00532_));
 BUF_X4 clkbuf_level_0_1_19__00532_ (.A(clknet_2_0__leaf__00532_),
    .Z(clknet_level_0_1_19__00532_));
 BUF_X4 clkbuf_level_1_1_110__00532_ (.A(clknet_level_0_1_19__00532_),
    .Z(clknet_level_1_1_110__00532_));
 BUF_X4 clkbuf_level_2_1_111__00532_ (.A(clknet_level_1_1_110__00532_),
    .Z(clknet_level_2_1_111__00532_));
 BUF_X4 clkbuf_level_3_1_112__00532_ (.A(clknet_level_2_1_111__00532_),
    .Z(clknet_level_3_1_112__00532_));
 BUF_X4 clkbuf_level_4_1_113__00532_ (.A(clknet_level_3_1_112__00532_),
    .Z(clknet_level_4_1_113__00532_));
 BUF_X4 clkbuf_level_5_1_114__00532_ (.A(clknet_level_4_1_113__00532_),
    .Z(clknet_level_5_1_114__00532_));
 BUF_X4 clkbuf_level_0_1_2111__00532_ (.A(clknet_2_1__leaf__00532_),
    .Z(clknet_level_0_1_2111__00532_));
 BUF_X4 clkbuf_level_1_1_2112__00532_ (.A(clknet_level_0_1_2111__00532_),
    .Z(clknet_level_1_1_2112__00532_));
 BUF_X4 clkbuf_level_2_1_2113__00532_ (.A(clknet_level_1_1_2112__00532_),
    .Z(clknet_level_2_1_2113__00532_));
 BUF_X4 clkbuf_level_3_1_2114__00532_ (.A(clknet_level_2_1_2113__00532_),
    .Z(clknet_level_3_1_2114__00532_));
 BUF_X4 clkbuf_level_4_1_2115__00532_ (.A(clknet_level_3_1_2114__00532_),
    .Z(clknet_level_4_1_2115__00532_));
 BUF_X4 clkbuf_level_5_1_2116__00532_ (.A(clknet_level_4_1_2115__00532_),
    .Z(clknet_level_5_1_2116__00532_));
 BUF_X4 clkbuf_level_0_1_3213__00532_ (.A(clknet_2_2__leaf__00532_),
    .Z(clknet_level_0_1_3213__00532_));
 BUF_X4 clkbuf_level_1_1_3214__00532_ (.A(clknet_level_0_1_3213__00532_),
    .Z(clknet_level_1_1_3214__00532_));
 BUF_X4 clkbuf_level_2_1_3215__00532_ (.A(clknet_level_1_1_3214__00532_),
    .Z(clknet_level_2_1_3215__00532_));
 BUF_X4 clkbuf_level_3_1_3216__00532_ (.A(clknet_level_2_1_3215__00532_),
    .Z(clknet_level_3_1_3216__00532_));
 BUF_X4 clkbuf_level_4_1_3217__00532_ (.A(clknet_level_3_1_3216__00532_),
    .Z(clknet_level_4_1_3217__00532_));
 BUF_X4 clkbuf_level_5_1_3218__00532_ (.A(clknet_level_4_1_3217__00532_),
    .Z(clknet_level_5_1_3218__00532_));
 BUF_X4 clkbuf_level_0_1_4315__00532_ (.A(clknet_2_3__leaf__00532_),
    .Z(clknet_level_0_1_4315__00532_));
 BUF_X4 clkbuf_level_1_1_4316__00532_ (.A(clknet_level_0_1_4315__00532_),
    .Z(clknet_level_1_1_4316__00532_));
 BUF_X4 clkbuf_level_2_1_4317__00532_ (.A(clknet_level_1_1_4316__00532_),
    .Z(clknet_level_2_1_4317__00532_));
 BUF_X4 clkbuf_level_3_1_4318__00532_ (.A(clknet_level_2_1_4317__00532_),
    .Z(clknet_level_3_1_4318__00532_));
 BUF_X4 clkbuf_level_4_1_4319__00532_ (.A(clknet_level_3_1_4318__00532_),
    .Z(clknet_level_4_1_4319__00532_));
 BUF_X4 clkbuf_level_5_1_4320__00532_ (.A(clknet_level_4_1_4319__00532_),
    .Z(clknet_level_5_1_4320__00532_));
 BUF_X4 clkbuf_0__00534_ (.A(_00534_),
    .Z(clknet_0__00534_));
 BUF_X4 clkbuf_3_0__f__00534_ (.A(clknet_0__00534_),
    .Z(clknet_3_0__leaf__00534_));
 BUF_X4 clkbuf_3_1__f__00534_ (.A(clknet_0__00534_),
    .Z(clknet_3_1__leaf__00534_));
 BUF_X4 clkbuf_3_2__f__00534_ (.A(clknet_0__00534_),
    .Z(clknet_3_2__leaf__00534_));
 BUF_X4 clkbuf_3_3__f__00534_ (.A(clknet_0__00534_),
    .Z(clknet_3_3__leaf__00534_));
 BUF_X4 clkbuf_3_4__f__00534_ (.A(clknet_0__00534_),
    .Z(clknet_3_4__leaf__00534_));
 BUF_X4 clkbuf_3_5__f__00534_ (.A(clknet_0__00534_),
    .Z(clknet_3_5__leaf__00534_));
 BUF_X4 clkbuf_3_6__f__00534_ (.A(clknet_0__00534_),
    .Z(clknet_3_6__leaf__00534_));
 BUF_X4 clkbuf_3_7__f__00534_ (.A(clknet_0__00534_),
    .Z(clknet_3_7__leaf__00534_));
 BUF_X4 clkbuf_level_0_1_1219__00534_ (.A(clknet_3_0__leaf__00534_),
    .Z(clknet_level_0_1_1219__00534_));
 BUF_X4 clkbuf_level_1_1_1220__00534_ (.A(clknet_level_0_1_1219__00534_),
    .Z(clknet_level_1_1_1220__00534_));
 BUF_X4 clkbuf_level_2_1_1221__00534_ (.A(clknet_level_1_1_1220__00534_),
    .Z(clknet_level_2_1_1221__00534_));
 BUF_X4 clkbuf_level_0_1_2222__00534_ (.A(clknet_3_1__leaf__00534_),
    .Z(clknet_level_0_1_2222__00534_));
 BUF_X4 clkbuf_level_1_1_2223__00534_ (.A(clknet_level_0_1_2222__00534_),
    .Z(clknet_level_1_1_2223__00534_));
 BUF_X4 clkbuf_level_2_1_2224__00534_ (.A(clknet_level_1_1_2223__00534_),
    .Z(clknet_level_2_1_2224__00534_));
 BUF_X4 clkbuf_level_0_1_3225__00534_ (.A(clknet_3_2__leaf__00534_),
    .Z(clknet_level_0_1_3225__00534_));
 BUF_X4 clkbuf_level_1_1_3226__00534_ (.A(clknet_level_0_1_3225__00534_),
    .Z(clknet_level_1_1_3226__00534_));
 BUF_X4 clkbuf_level_2_1_3227__00534_ (.A(clknet_level_1_1_3226__00534_),
    .Z(clknet_level_2_1_3227__00534_));
 BUF_X4 clkbuf_level_0_1_4228__00534_ (.A(clknet_3_3__leaf__00534_),
    .Z(clknet_level_0_1_4228__00534_));
 BUF_X4 clkbuf_level_1_1_4229__00534_ (.A(clknet_level_0_1_4228__00534_),
    .Z(clknet_level_1_1_4229__00534_));
 BUF_X4 clkbuf_level_2_1_4230__00534_ (.A(clknet_level_1_1_4229__00534_),
    .Z(clknet_level_2_1_4230__00534_));
 BUF_X4 clkbuf_level_0_1_5231__00534_ (.A(clknet_3_4__leaf__00534_),
    .Z(clknet_level_0_1_5231__00534_));
 BUF_X4 clkbuf_level_1_1_5232__00534_ (.A(clknet_level_0_1_5231__00534_),
    .Z(clknet_level_1_1_5232__00534_));
 BUF_X4 clkbuf_level_2_1_5233__00534_ (.A(clknet_level_1_1_5232__00534_),
    .Z(clknet_level_2_1_5233__00534_));
 BUF_X4 clkbuf_level_0_1_6234__00534_ (.A(clknet_3_5__leaf__00534_),
    .Z(clknet_level_0_1_6234__00534_));
 BUF_X4 clkbuf_level_1_1_6235__00534_ (.A(clknet_level_0_1_6234__00534_),
    .Z(clknet_level_1_1_6235__00534_));
 BUF_X4 clkbuf_level_2_1_6236__00534_ (.A(clknet_level_1_1_6235__00534_),
    .Z(clknet_level_2_1_6236__00534_));
 BUF_X4 clkbuf_level_0_1_7237__00534_ (.A(clknet_3_6__leaf__00534_),
    .Z(clknet_level_0_1_7237__00534_));
 BUF_X4 clkbuf_level_1_1_7238__00534_ (.A(clknet_level_0_1_7237__00534_),
    .Z(clknet_level_1_1_7238__00534_));
 BUF_X4 clkbuf_level_2_1_7239__00534_ (.A(clknet_level_1_1_7238__00534_),
    .Z(clknet_level_2_1_7239__00534_));
 BUF_X4 clkbuf_level_0_1_8240__00534_ (.A(clknet_3_7__leaf__00534_),
    .Z(clknet_level_0_1_8240__00534_));
 BUF_X4 clkbuf_level_1_1_8241__00534_ (.A(clknet_level_0_1_8240__00534_),
    .Z(clknet_level_1_1_8241__00534_));
 BUF_X4 clkbuf_level_2_1_8242__00534_ (.A(clknet_level_1_1_8241__00534_),
    .Z(clknet_level_2_1_8242__00534_));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__15.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ));
 BUF_X4 clkbuf_0__00537_ (.A(_00537_),
    .Z(clknet_0__00537_));
 BUF_X4 clkbuf_3_0__f__00537_ (.A(clknet_0__00537_),
    .Z(clknet_3_0__leaf__00537_));
 BUF_X4 clkbuf_3_1__f__00537_ (.A(clknet_0__00537_),
    .Z(clknet_3_1__leaf__00537_));
 BUF_X4 clkbuf_3_2__f__00537_ (.A(clknet_0__00537_),
    .Z(clknet_3_2__leaf__00537_));
 BUF_X4 clkbuf_3_3__f__00537_ (.A(clknet_0__00537_),
    .Z(clknet_3_3__leaf__00537_));
 BUF_X4 clkbuf_3_4__f__00537_ (.A(clknet_0__00537_),
    .Z(clknet_3_4__leaf__00537_));
 BUF_X4 clkbuf_3_5__f__00537_ (.A(clknet_0__00537_),
    .Z(clknet_3_5__leaf__00537_));
 BUF_X4 clkbuf_3_6__f__00537_ (.A(clknet_0__00537_),
    .Z(clknet_3_6__leaf__00537_));
 BUF_X4 clkbuf_3_7__f__00537_ (.A(clknet_0__00537_),
    .Z(clknet_3_7__leaf__00537_));
 BUF_X4 clkbuf_level_0_1_1117__00537_ (.A(clknet_3_0__leaf__00537_),
    .Z(clknet_level_0_1_1117__00537_));
 BUF_X4 clkbuf_level_1_1_1118__00537_ (.A(clknet_level_0_1_1117__00537_),
    .Z(clknet_level_1_1_1118__00537_));
 BUF_X4 clkbuf_level_2_1_1119__00537_ (.A(clknet_level_1_1_1118__00537_),
    .Z(clknet_level_2_1_1119__00537_));
 BUF_X4 clkbuf_level_0_1_2120__00537_ (.A(clknet_3_1__leaf__00537_),
    .Z(clknet_level_0_1_2120__00537_));
 BUF_X4 clkbuf_level_1_1_2121__00537_ (.A(clknet_level_0_1_2120__00537_),
    .Z(clknet_level_1_1_2121__00537_));
 BUF_X4 clkbuf_level_2_1_2122__00537_ (.A(clknet_level_1_1_2121__00537_),
    .Z(clknet_level_2_1_2122__00537_));
 BUF_X4 clkbuf_level_0_1_3123__00537_ (.A(clknet_3_2__leaf__00537_),
    .Z(clknet_level_0_1_3123__00537_));
 BUF_X4 clkbuf_level_1_1_3124__00537_ (.A(clknet_level_0_1_3123__00537_),
    .Z(clknet_level_1_1_3124__00537_));
 BUF_X4 clkbuf_level_2_1_3125__00537_ (.A(clknet_level_1_1_3124__00537_),
    .Z(clknet_level_2_1_3125__00537_));
 BUF_X4 clkbuf_level_0_1_4126__00537_ (.A(clknet_3_3__leaf__00537_),
    .Z(clknet_level_0_1_4126__00537_));
 BUF_X4 clkbuf_level_1_1_4127__00537_ (.A(clknet_level_0_1_4126__00537_),
    .Z(clknet_level_1_1_4127__00537_));
 BUF_X4 clkbuf_level_2_1_4128__00537_ (.A(clknet_level_1_1_4127__00537_),
    .Z(clknet_level_2_1_4128__00537_));
 BUF_X4 clkbuf_level_0_1_5129__00537_ (.A(clknet_3_4__leaf__00537_),
    .Z(clknet_level_0_1_5129__00537_));
 BUF_X4 clkbuf_level_1_1_5130__00537_ (.A(clknet_level_0_1_5129__00537_),
    .Z(clknet_level_1_1_5130__00537_));
 BUF_X4 clkbuf_level_2_1_5131__00537_ (.A(clknet_level_1_1_5130__00537_),
    .Z(clknet_level_2_1_5131__00537_));
 BUF_X4 clkbuf_level_0_1_6132__00537_ (.A(clknet_3_5__leaf__00537_),
    .Z(clknet_level_0_1_6132__00537_));
 BUF_X4 clkbuf_level_1_1_6133__00537_ (.A(clknet_level_0_1_6132__00537_),
    .Z(clknet_level_1_1_6133__00537_));
 BUF_X4 clkbuf_level_2_1_6134__00537_ (.A(clknet_level_1_1_6133__00537_),
    .Z(clknet_level_2_1_6134__00537_));
 BUF_X4 clkbuf_level_0_1_7135__00537_ (.A(clknet_3_6__leaf__00537_),
    .Z(clknet_level_0_1_7135__00537_));
 BUF_X4 clkbuf_level_1_1_7136__00537_ (.A(clknet_level_0_1_7135__00537_),
    .Z(clknet_level_1_1_7136__00537_));
 BUF_X4 clkbuf_level_2_1_7137__00537_ (.A(clknet_level_1_1_7136__00537_),
    .Z(clknet_level_2_1_7137__00537_));
 BUF_X4 clkbuf_level_0_1_8138__00537_ (.A(clknet_3_7__leaf__00537_),
    .Z(clknet_level_0_1_8138__00537_));
 BUF_X4 clkbuf_level_1_1_8139__00537_ (.A(clknet_level_0_1_8138__00537_),
    .Z(clknet_level_1_1_8139__00537_));
 BUF_X4 clkbuf_level_2_1_8140__00537_ (.A(clknet_level_1_1_8139__00537_),
    .Z(clknet_level_2_1_8140__00537_));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__14.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ));
 BUF_X4 clkbuf_0__00540_ (.A(_00540_),
    .Z(clknet_0__00540_));
 BUF_X4 clkbuf_3_0__f__00540_ (.A(clknet_0__00540_),
    .Z(clknet_3_0__leaf__00540_));
 BUF_X4 clkbuf_3_1__f__00540_ (.A(clknet_0__00540_),
    .Z(clknet_3_1__leaf__00540_));
 BUF_X4 clkbuf_3_2__f__00540_ (.A(clknet_0__00540_),
    .Z(clknet_3_2__leaf__00540_));
 BUF_X4 clkbuf_3_3__f__00540_ (.A(clknet_0__00540_),
    .Z(clknet_3_3__leaf__00540_));
 BUF_X4 clkbuf_3_4__f__00540_ (.A(clknet_0__00540_),
    .Z(clknet_3_4__leaf__00540_));
 BUF_X4 clkbuf_3_5__f__00540_ (.A(clknet_0__00540_),
    .Z(clknet_3_5__leaf__00540_));
 BUF_X4 clkbuf_3_6__f__00540_ (.A(clknet_0__00540_),
    .Z(clknet_3_6__leaf__00540_));
 BUF_X4 clkbuf_3_7__f__00540_ (.A(clknet_0__00540_),
    .Z(clknet_3_7__leaf__00540_));
 BUF_X4 clkbuf_level_0_1_1321__00540_ (.A(clknet_3_0__leaf__00540_),
    .Z(clknet_level_0_1_1321__00540_));
 BUF_X4 clkbuf_level_1_1_1322__00540_ (.A(clknet_level_0_1_1321__00540_),
    .Z(clknet_level_1_1_1322__00540_));
 BUF_X4 clkbuf_level_2_1_1323__00540_ (.A(clknet_level_1_1_1322__00540_),
    .Z(clknet_level_2_1_1323__00540_));
 BUF_X4 clkbuf_level_0_1_2324__00540_ (.A(clknet_3_1__leaf__00540_),
    .Z(clknet_level_0_1_2324__00540_));
 BUF_X4 clkbuf_level_1_1_2325__00540_ (.A(clknet_level_0_1_2324__00540_),
    .Z(clknet_level_1_1_2325__00540_));
 BUF_X4 clkbuf_level_2_1_2326__00540_ (.A(clknet_level_1_1_2325__00540_),
    .Z(clknet_level_2_1_2326__00540_));
 BUF_X4 clkbuf_level_0_1_3327__00540_ (.A(clknet_3_2__leaf__00540_),
    .Z(clknet_level_0_1_3327__00540_));
 BUF_X4 clkbuf_level_1_1_3328__00540_ (.A(clknet_level_0_1_3327__00540_),
    .Z(clknet_level_1_1_3328__00540_));
 BUF_X4 clkbuf_level_2_1_3329__00540_ (.A(clknet_level_1_1_3328__00540_),
    .Z(clknet_level_2_1_3329__00540_));
 BUF_X4 clkbuf_level_0_1_4330__00540_ (.A(clknet_3_3__leaf__00540_),
    .Z(clknet_level_0_1_4330__00540_));
 BUF_X4 clkbuf_level_1_1_4331__00540_ (.A(clknet_level_0_1_4330__00540_),
    .Z(clknet_level_1_1_4331__00540_));
 BUF_X4 clkbuf_level_2_1_4332__00540_ (.A(clknet_level_1_1_4331__00540_),
    .Z(clknet_level_2_1_4332__00540_));
 BUF_X4 clkbuf_level_0_1_5333__00540_ (.A(clknet_3_4__leaf__00540_),
    .Z(clknet_level_0_1_5333__00540_));
 BUF_X4 clkbuf_level_1_1_5334__00540_ (.A(clknet_level_0_1_5333__00540_),
    .Z(clknet_level_1_1_5334__00540_));
 BUF_X4 clkbuf_level_2_1_5335__00540_ (.A(clknet_level_1_1_5334__00540_),
    .Z(clknet_level_2_1_5335__00540_));
 BUF_X4 clkbuf_level_0_1_6336__00540_ (.A(clknet_3_5__leaf__00540_),
    .Z(clknet_level_0_1_6336__00540_));
 BUF_X4 clkbuf_level_1_1_6337__00540_ (.A(clknet_level_0_1_6336__00540_),
    .Z(clknet_level_1_1_6337__00540_));
 BUF_X4 clkbuf_level_2_1_6338__00540_ (.A(clknet_level_1_1_6337__00540_),
    .Z(clknet_level_2_1_6338__00540_));
 BUF_X4 clkbuf_level_0_1_7339__00540_ (.A(clknet_3_6__leaf__00540_),
    .Z(clknet_level_0_1_7339__00540_));
 BUF_X4 clkbuf_level_1_1_7340__00540_ (.A(clknet_level_0_1_7339__00540_),
    .Z(clknet_level_1_1_7340__00540_));
 BUF_X4 clkbuf_level_2_1_7341__00540_ (.A(clknet_level_1_1_7340__00540_),
    .Z(clknet_level_2_1_7341__00540_));
 BUF_X4 clkbuf_level_0_1_8342__00540_ (.A(clknet_3_7__leaf__00540_),
    .Z(clknet_level_0_1_8342__00540_));
 BUF_X4 clkbuf_level_1_1_8343__00540_ (.A(clknet_level_0_1_8342__00540_),
    .Z(clknet_level_1_1_8343__00540_));
 BUF_X4 clkbuf_level_2_1_8344__00540_ (.A(clknet_level_1_1_8343__00540_),
    .Z(clknet_level_2_1_8344__00540_));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__13.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ));
 BUF_X4 clkbuf_0__00543_ (.A(_00543_),
    .Z(clknet_0__00543_));
 BUF_X4 clkbuf_3_0__f__00543_ (.A(clknet_0__00543_),
    .Z(clknet_3_0__leaf__00543_));
 BUF_X4 clkbuf_3_1__f__00543_ (.A(clknet_0__00543_),
    .Z(clknet_3_1__leaf__00543_));
 BUF_X4 clkbuf_3_2__f__00543_ (.A(clknet_0__00543_),
    .Z(clknet_3_2__leaf__00543_));
 BUF_X4 clkbuf_3_3__f__00543_ (.A(clknet_0__00543_),
    .Z(clknet_3_3__leaf__00543_));
 BUF_X4 clkbuf_3_4__f__00543_ (.A(clknet_0__00543_),
    .Z(clknet_3_4__leaf__00543_));
 BUF_X4 clkbuf_3_5__f__00543_ (.A(clknet_0__00543_),
    .Z(clknet_3_5__leaf__00543_));
 BUF_X4 clkbuf_3_6__f__00543_ (.A(clknet_0__00543_),
    .Z(clknet_3_6__leaf__00543_));
 BUF_X4 clkbuf_3_7__f__00543_ (.A(clknet_0__00543_),
    .Z(clknet_3_7__leaf__00543_));
 BUF_X4 clkbuf_level_0_1_1141__00543_ (.A(clknet_3_0__leaf__00543_),
    .Z(clknet_level_0_1_1141__00543_));
 BUF_X4 clkbuf_level_1_1_1142__00543_ (.A(clknet_level_0_1_1141__00543_),
    .Z(clknet_level_1_1_1142__00543_));
 BUF_X4 clkbuf_level_2_1_1143__00543_ (.A(clknet_level_1_1_1142__00543_),
    .Z(clknet_level_2_1_1143__00543_));
 BUF_X4 clkbuf_level_0_1_2144__00543_ (.A(clknet_3_1__leaf__00543_),
    .Z(clknet_level_0_1_2144__00543_));
 BUF_X4 clkbuf_level_1_1_2145__00543_ (.A(clknet_level_0_1_2144__00543_),
    .Z(clknet_level_1_1_2145__00543_));
 BUF_X4 clkbuf_level_2_1_2146__00543_ (.A(clknet_level_1_1_2145__00543_),
    .Z(clknet_level_2_1_2146__00543_));
 BUF_X4 clkbuf_level_0_1_3147__00543_ (.A(clknet_3_2__leaf__00543_),
    .Z(clknet_level_0_1_3147__00543_));
 BUF_X4 clkbuf_level_1_1_3148__00543_ (.A(clknet_level_0_1_3147__00543_),
    .Z(clknet_level_1_1_3148__00543_));
 BUF_X4 clkbuf_level_2_1_3149__00543_ (.A(clknet_level_1_1_3148__00543_),
    .Z(clknet_level_2_1_3149__00543_));
 BUF_X4 clkbuf_level_0_1_4150__00543_ (.A(clknet_3_3__leaf__00543_),
    .Z(clknet_level_0_1_4150__00543_));
 BUF_X4 clkbuf_level_1_1_4151__00543_ (.A(clknet_level_0_1_4150__00543_),
    .Z(clknet_level_1_1_4151__00543_));
 BUF_X4 clkbuf_level_2_1_4152__00543_ (.A(clknet_level_1_1_4151__00543_),
    .Z(clknet_level_2_1_4152__00543_));
 BUF_X4 clkbuf_level_0_1_5153__00543_ (.A(clknet_3_4__leaf__00543_),
    .Z(clknet_level_0_1_5153__00543_));
 BUF_X4 clkbuf_level_1_1_5154__00543_ (.A(clknet_level_0_1_5153__00543_),
    .Z(clknet_level_1_1_5154__00543_));
 BUF_X4 clkbuf_level_2_1_5155__00543_ (.A(clknet_level_1_1_5154__00543_),
    .Z(clknet_level_2_1_5155__00543_));
 BUF_X4 clkbuf_level_0_1_6156__00543_ (.A(clknet_3_5__leaf__00543_),
    .Z(clknet_level_0_1_6156__00543_));
 BUF_X4 clkbuf_level_1_1_6157__00543_ (.A(clknet_level_0_1_6156__00543_),
    .Z(clknet_level_1_1_6157__00543_));
 BUF_X4 clkbuf_level_2_1_6158__00543_ (.A(clknet_level_1_1_6157__00543_),
    .Z(clknet_level_2_1_6158__00543_));
 BUF_X4 clkbuf_level_0_1_7159__00543_ (.A(clknet_3_6__leaf__00543_),
    .Z(clknet_level_0_1_7159__00543_));
 BUF_X4 clkbuf_level_1_1_7160__00543_ (.A(clknet_level_0_1_7159__00543_),
    .Z(clknet_level_1_1_7160__00543_));
 BUF_X4 clkbuf_level_2_1_7161__00543_ (.A(clknet_level_1_1_7160__00543_),
    .Z(clknet_level_2_1_7161__00543_));
 BUF_X4 clkbuf_level_0_1_8162__00543_ (.A(clknet_3_7__leaf__00543_),
    .Z(clknet_level_0_1_8162__00543_));
 BUF_X4 clkbuf_level_1_1_8163__00543_ (.A(clknet_level_0_1_8162__00543_),
    .Z(clknet_level_1_1_8163__00543_));
 BUF_X4 clkbuf_level_2_1_8164__00543_ (.A(clknet_level_1_1_8163__00543_),
    .Z(clknet_level_2_1_8164__00543_));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__12.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ));
 BUF_X4 clkbuf_0__00546_ (.A(_00546_),
    .Z(clknet_0__00546_));
 BUF_X4 clkbuf_3_0__f__00546_ (.A(clknet_0__00546_),
    .Z(clknet_3_0__leaf__00546_));
 BUF_X4 clkbuf_3_1__f__00546_ (.A(clknet_0__00546_),
    .Z(clknet_3_1__leaf__00546_));
 BUF_X4 clkbuf_3_2__f__00546_ (.A(clknet_0__00546_),
    .Z(clknet_3_2__leaf__00546_));
 BUF_X4 clkbuf_3_3__f__00546_ (.A(clknet_0__00546_),
    .Z(clknet_3_3__leaf__00546_));
 BUF_X4 clkbuf_3_4__f__00546_ (.A(clknet_0__00546_),
    .Z(clknet_3_4__leaf__00546_));
 BUF_X4 clkbuf_3_5__f__00546_ (.A(clknet_0__00546_),
    .Z(clknet_3_5__leaf__00546_));
 BUF_X4 clkbuf_3_6__f__00546_ (.A(clknet_0__00546_),
    .Z(clknet_3_6__leaf__00546_));
 BUF_X4 clkbuf_3_7__f__00546_ (.A(clknet_0__00546_),
    .Z(clknet_3_7__leaf__00546_));
 BUF_X4 clkbuf_level_0_1_1345__00546_ (.A(clknet_3_0__leaf__00546_),
    .Z(clknet_level_0_1_1345__00546_));
 BUF_X4 clkbuf_level_1_1_1346__00546_ (.A(clknet_level_0_1_1345__00546_),
    .Z(clknet_level_1_1_1346__00546_));
 BUF_X4 clkbuf_level_2_1_1347__00546_ (.A(clknet_level_1_1_1346__00546_),
    .Z(clknet_level_2_1_1347__00546_));
 BUF_X4 clkbuf_level_0_1_2348__00546_ (.A(clknet_3_1__leaf__00546_),
    .Z(clknet_level_0_1_2348__00546_));
 BUF_X4 clkbuf_level_1_1_2349__00546_ (.A(clknet_level_0_1_2348__00546_),
    .Z(clknet_level_1_1_2349__00546_));
 BUF_X4 clkbuf_level_2_1_2350__00546_ (.A(clknet_level_1_1_2349__00546_),
    .Z(clknet_level_2_1_2350__00546_));
 BUF_X4 clkbuf_level_0_1_3351__00546_ (.A(clknet_3_2__leaf__00546_),
    .Z(clknet_level_0_1_3351__00546_));
 BUF_X4 clkbuf_level_1_1_3352__00546_ (.A(clknet_level_0_1_3351__00546_),
    .Z(clknet_level_1_1_3352__00546_));
 BUF_X4 clkbuf_level_2_1_3353__00546_ (.A(clknet_level_1_1_3352__00546_),
    .Z(clknet_level_2_1_3353__00546_));
 BUF_X4 clkbuf_level_0_1_4354__00546_ (.A(clknet_3_3__leaf__00546_),
    .Z(clknet_level_0_1_4354__00546_));
 BUF_X4 clkbuf_level_1_1_4355__00546_ (.A(clknet_level_0_1_4354__00546_),
    .Z(clknet_level_1_1_4355__00546_));
 BUF_X4 clkbuf_level_2_1_4356__00546_ (.A(clknet_level_1_1_4355__00546_),
    .Z(clknet_level_2_1_4356__00546_));
 BUF_X4 clkbuf_level_0_1_5357__00546_ (.A(clknet_3_4__leaf__00546_),
    .Z(clknet_level_0_1_5357__00546_));
 BUF_X4 clkbuf_level_1_1_5358__00546_ (.A(clknet_level_0_1_5357__00546_),
    .Z(clknet_level_1_1_5358__00546_));
 BUF_X4 clkbuf_level_2_1_5359__00546_ (.A(clknet_level_1_1_5358__00546_),
    .Z(clknet_level_2_1_5359__00546_));
 BUF_X4 clkbuf_level_0_1_6360__00546_ (.A(clknet_3_5__leaf__00546_),
    .Z(clknet_level_0_1_6360__00546_));
 BUF_X4 clkbuf_level_1_1_6361__00546_ (.A(clknet_level_0_1_6360__00546_),
    .Z(clknet_level_1_1_6361__00546_));
 BUF_X4 clkbuf_level_2_1_6362__00546_ (.A(clknet_level_1_1_6361__00546_),
    .Z(clknet_level_2_1_6362__00546_));
 BUF_X4 clkbuf_level_0_1_7363__00546_ (.A(clknet_3_6__leaf__00546_),
    .Z(clknet_level_0_1_7363__00546_));
 BUF_X4 clkbuf_level_1_1_7364__00546_ (.A(clknet_level_0_1_7363__00546_),
    .Z(clknet_level_1_1_7364__00546_));
 BUF_X4 clkbuf_level_2_1_7365__00546_ (.A(clknet_level_1_1_7364__00546_),
    .Z(clknet_level_2_1_7365__00546_));
 BUF_X4 clkbuf_level_0_1_8366__00546_ (.A(clknet_3_7__leaf__00546_),
    .Z(clknet_level_0_1_8366__00546_));
 BUF_X4 clkbuf_level_1_1_8367__00546_ (.A(clknet_level_0_1_8366__00546_),
    .Z(clknet_level_1_1_8367__00546_));
 BUF_X4 clkbuf_level_2_1_8368__00546_ (.A(clknet_level_1_1_8367__00546_),
    .Z(clknet_level_2_1_8368__00546_));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__11.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ));
 BUF_X4 clkbuf_0__00549_ (.A(_00549_),
    .Z(clknet_0__00549_));
 BUF_X4 clkbuf_3_0__f__00549_ (.A(clknet_0__00549_),
    .Z(clknet_3_0__leaf__00549_));
 BUF_X4 clkbuf_3_1__f__00549_ (.A(clknet_0__00549_),
    .Z(clknet_3_1__leaf__00549_));
 BUF_X4 clkbuf_3_2__f__00549_ (.A(clknet_0__00549_),
    .Z(clknet_3_2__leaf__00549_));
 BUF_X4 clkbuf_3_3__f__00549_ (.A(clknet_0__00549_),
    .Z(clknet_3_3__leaf__00549_));
 BUF_X4 clkbuf_3_4__f__00549_ (.A(clknet_0__00549_),
    .Z(clknet_3_4__leaf__00549_));
 BUF_X4 clkbuf_3_5__f__00549_ (.A(clknet_0__00549_),
    .Z(clknet_3_5__leaf__00549_));
 BUF_X4 clkbuf_3_6__f__00549_ (.A(clknet_0__00549_),
    .Z(clknet_3_6__leaf__00549_));
 BUF_X4 clkbuf_3_7__f__00549_ (.A(clknet_0__00549_),
    .Z(clknet_3_7__leaf__00549_));
 BUF_X4 clkbuf_level_0_1_115__00549_ (.A(clknet_3_0__leaf__00549_),
    .Z(clknet_level_0_1_115__00549_));
 BUF_X4 clkbuf_level_1_1_116__00549_ (.A(clknet_level_0_1_115__00549_),
    .Z(clknet_level_1_1_116__00549_));
 BUF_X4 clkbuf_level_2_1_117__00549_ (.A(clknet_level_1_1_116__00549_),
    .Z(clknet_level_2_1_117__00549_));
 BUF_X4 clkbuf_level_0_1_218__00549_ (.A(clknet_3_1__leaf__00549_),
    .Z(clknet_level_0_1_218__00549_));
 BUF_X4 clkbuf_level_1_1_219__00549_ (.A(clknet_level_0_1_218__00549_),
    .Z(clknet_level_1_1_219__00549_));
 BUF_X4 clkbuf_level_2_1_220__00549_ (.A(clknet_level_1_1_219__00549_),
    .Z(clknet_level_2_1_220__00549_));
 BUF_X4 clkbuf_level_0_1_321__00549_ (.A(clknet_3_2__leaf__00549_),
    .Z(clknet_level_0_1_321__00549_));
 BUF_X4 clkbuf_level_1_1_322__00549_ (.A(clknet_level_0_1_321__00549_),
    .Z(clknet_level_1_1_322__00549_));
 BUF_X4 clkbuf_level_2_1_323__00549_ (.A(clknet_level_1_1_322__00549_),
    .Z(clknet_level_2_1_323__00549_));
 BUF_X4 clkbuf_level_0_1_424__00549_ (.A(clknet_3_3__leaf__00549_),
    .Z(clknet_level_0_1_424__00549_));
 BUF_X4 clkbuf_level_1_1_425__00549_ (.A(clknet_level_0_1_424__00549_),
    .Z(clknet_level_1_1_425__00549_));
 BUF_X4 clkbuf_level_2_1_426__00549_ (.A(clknet_level_1_1_425__00549_),
    .Z(clknet_level_2_1_426__00549_));
 BUF_X4 clkbuf_level_0_1_527__00549_ (.A(clknet_3_4__leaf__00549_),
    .Z(clknet_level_0_1_527__00549_));
 BUF_X4 clkbuf_level_1_1_528__00549_ (.A(clknet_level_0_1_527__00549_),
    .Z(clknet_level_1_1_528__00549_));
 BUF_X4 clkbuf_level_2_1_529__00549_ (.A(clknet_level_1_1_528__00549_),
    .Z(clknet_level_2_1_529__00549_));
 BUF_X4 clkbuf_level_0_1_630__00549_ (.A(clknet_3_5__leaf__00549_),
    .Z(clknet_level_0_1_630__00549_));
 BUF_X4 clkbuf_level_1_1_631__00549_ (.A(clknet_level_0_1_630__00549_),
    .Z(clknet_level_1_1_631__00549_));
 BUF_X4 clkbuf_level_2_1_632__00549_ (.A(clknet_level_1_1_631__00549_),
    .Z(clknet_level_2_1_632__00549_));
 BUF_X4 clkbuf_level_0_1_733__00549_ (.A(clknet_3_6__leaf__00549_),
    .Z(clknet_level_0_1_733__00549_));
 BUF_X4 clkbuf_level_1_1_734__00549_ (.A(clknet_level_0_1_733__00549_),
    .Z(clknet_level_1_1_734__00549_));
 BUF_X4 clkbuf_level_2_1_735__00549_ (.A(clknet_level_1_1_734__00549_),
    .Z(clknet_level_2_1_735__00549_));
 BUF_X4 clkbuf_level_0_1_836__00549_ (.A(clknet_3_7__leaf__00549_),
    .Z(clknet_level_0_1_836__00549_));
 BUF_X4 clkbuf_level_1_1_837__00549_ (.A(clknet_level_0_1_836__00549_),
    .Z(clknet_level_1_1_837__00549_));
 BUF_X4 clkbuf_level_2_1_838__00549_ (.A(clknet_level_1_1_837__00549_),
    .Z(clknet_level_2_1_838__00549_));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__10.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ));
 BUF_X4 clkbuf_0__00552_ (.A(_00552_),
    .Z(clknet_0__00552_));
 BUF_X4 clkbuf_3_0__f__00552_ (.A(clknet_0__00552_),
    .Z(clknet_3_0__leaf__00552_));
 BUF_X4 clkbuf_3_1__f__00552_ (.A(clknet_0__00552_),
    .Z(clknet_3_1__leaf__00552_));
 BUF_X4 clkbuf_3_2__f__00552_ (.A(clknet_0__00552_),
    .Z(clknet_3_2__leaf__00552_));
 BUF_X4 clkbuf_3_3__f__00552_ (.A(clknet_0__00552_),
    .Z(clknet_3_3__leaf__00552_));
 BUF_X4 clkbuf_3_4__f__00552_ (.A(clknet_0__00552_),
    .Z(clknet_3_4__leaf__00552_));
 BUF_X4 clkbuf_3_5__f__00552_ (.A(clknet_0__00552_),
    .Z(clknet_3_5__leaf__00552_));
 BUF_X4 clkbuf_3_6__f__00552_ (.A(clknet_0__00552_),
    .Z(clknet_3_6__leaf__00552_));
 BUF_X4 clkbuf_3_7__f__00552_ (.A(clknet_0__00552_),
    .Z(clknet_3_7__leaf__00552_));
 BUF_X4 clkbuf_level_0_1_1165__00552_ (.A(clknet_3_0__leaf__00552_),
    .Z(clknet_level_0_1_1165__00552_));
 BUF_X4 clkbuf_level_1_1_1166__00552_ (.A(clknet_level_0_1_1165__00552_),
    .Z(clknet_level_1_1_1166__00552_));
 BUF_X4 clkbuf_level_2_1_1167__00552_ (.A(clknet_level_1_1_1166__00552_),
    .Z(clknet_level_2_1_1167__00552_));
 BUF_X4 clkbuf_level_0_1_2168__00552_ (.A(clknet_3_1__leaf__00552_),
    .Z(clknet_level_0_1_2168__00552_));
 BUF_X4 clkbuf_level_1_1_2169__00552_ (.A(clknet_level_0_1_2168__00552_),
    .Z(clknet_level_1_1_2169__00552_));
 BUF_X4 clkbuf_level_2_1_2170__00552_ (.A(clknet_level_1_1_2169__00552_),
    .Z(clknet_level_2_1_2170__00552_));
 BUF_X4 clkbuf_level_0_1_3171__00552_ (.A(clknet_3_2__leaf__00552_),
    .Z(clknet_level_0_1_3171__00552_));
 BUF_X4 clkbuf_level_1_1_3172__00552_ (.A(clknet_level_0_1_3171__00552_),
    .Z(clknet_level_1_1_3172__00552_));
 BUF_X4 clkbuf_level_2_1_3173__00552_ (.A(clknet_level_1_1_3172__00552_),
    .Z(clknet_level_2_1_3173__00552_));
 BUF_X4 clkbuf_level_0_1_4174__00552_ (.A(clknet_3_3__leaf__00552_),
    .Z(clknet_level_0_1_4174__00552_));
 BUF_X4 clkbuf_level_1_1_4175__00552_ (.A(clknet_level_0_1_4174__00552_),
    .Z(clknet_level_1_1_4175__00552_));
 BUF_X4 clkbuf_level_2_1_4176__00552_ (.A(clknet_level_1_1_4175__00552_),
    .Z(clknet_level_2_1_4176__00552_));
 BUF_X4 clkbuf_level_0_1_5177__00552_ (.A(clknet_3_4__leaf__00552_),
    .Z(clknet_level_0_1_5177__00552_));
 BUF_X4 clkbuf_level_1_1_5178__00552_ (.A(clknet_level_0_1_5177__00552_),
    .Z(clknet_level_1_1_5178__00552_));
 BUF_X4 clkbuf_level_2_1_5179__00552_ (.A(clknet_level_1_1_5178__00552_),
    .Z(clknet_level_2_1_5179__00552_));
 BUF_X4 clkbuf_level_0_1_6180__00552_ (.A(clknet_3_5__leaf__00552_),
    .Z(clknet_level_0_1_6180__00552_));
 BUF_X4 clkbuf_level_1_1_6181__00552_ (.A(clknet_level_0_1_6180__00552_),
    .Z(clknet_level_1_1_6181__00552_));
 BUF_X4 clkbuf_level_2_1_6182__00552_ (.A(clknet_level_1_1_6181__00552_),
    .Z(clknet_level_2_1_6182__00552_));
 BUF_X4 clkbuf_level_0_1_7183__00552_ (.A(clknet_3_6__leaf__00552_),
    .Z(clknet_level_0_1_7183__00552_));
 BUF_X4 clkbuf_level_1_1_7184__00552_ (.A(clknet_level_0_1_7183__00552_),
    .Z(clknet_level_1_1_7184__00552_));
 BUF_X4 clkbuf_level_2_1_7185__00552_ (.A(clknet_level_1_1_7184__00552_),
    .Z(clknet_level_2_1_7185__00552_));
 BUF_X4 clkbuf_level_0_1_8186__00552_ (.A(clknet_3_7__leaf__00552_),
    .Z(clknet_level_0_1_8186__00552_));
 BUF_X4 clkbuf_level_1_1_8187__00552_ (.A(clknet_level_0_1_8186__00552_),
    .Z(clknet_level_1_1_8187__00552_));
 BUF_X4 clkbuf_level_2_1_8188__00552_ (.A(clknet_level_1_1_8187__00552_),
    .Z(clknet_level_2_1_8188__00552_));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__9.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ));
 BUF_X4 clkbuf_0__00555_ (.A(_00555_),
    .Z(clknet_0__00555_));
 BUF_X4 clkbuf_3_0__f__00555_ (.A(clknet_0__00555_),
    .Z(clknet_3_0__leaf__00555_));
 BUF_X4 clkbuf_3_1__f__00555_ (.A(clknet_0__00555_),
    .Z(clknet_3_1__leaf__00555_));
 BUF_X4 clkbuf_3_2__f__00555_ (.A(clknet_0__00555_),
    .Z(clknet_3_2__leaf__00555_));
 BUF_X4 clkbuf_3_3__f__00555_ (.A(clknet_0__00555_),
    .Z(clknet_3_3__leaf__00555_));
 BUF_X4 clkbuf_3_4__f__00555_ (.A(clknet_0__00555_),
    .Z(clknet_3_4__leaf__00555_));
 BUF_X4 clkbuf_3_5__f__00555_ (.A(clknet_0__00555_),
    .Z(clknet_3_5__leaf__00555_));
 BUF_X4 clkbuf_3_6__f__00555_ (.A(clknet_0__00555_),
    .Z(clknet_3_6__leaf__00555_));
 BUF_X4 clkbuf_3_7__f__00555_ (.A(clknet_0__00555_),
    .Z(clknet_3_7__leaf__00555_));
 BUF_X4 clkbuf_level_0_1_139__00555_ (.A(clknet_3_0__leaf__00555_),
    .Z(clknet_level_0_1_139__00555_));
 BUF_X4 clkbuf_level_1_1_140__00555_ (.A(clknet_level_0_1_139__00555_),
    .Z(clknet_level_1_1_140__00555_));
 BUF_X4 clkbuf_level_2_1_141__00555_ (.A(clknet_level_1_1_140__00555_),
    .Z(clknet_level_2_1_141__00555_));
 BUF_X4 clkbuf_level_0_1_242__00555_ (.A(clknet_3_1__leaf__00555_),
    .Z(clknet_level_0_1_242__00555_));
 BUF_X4 clkbuf_level_1_1_243__00555_ (.A(clknet_level_0_1_242__00555_),
    .Z(clknet_level_1_1_243__00555_));
 BUF_X4 clkbuf_level_2_1_244__00555_ (.A(clknet_level_1_1_243__00555_),
    .Z(clknet_level_2_1_244__00555_));
 BUF_X4 clkbuf_level_0_1_345__00555_ (.A(clknet_3_2__leaf__00555_),
    .Z(clknet_level_0_1_345__00555_));
 BUF_X4 clkbuf_level_1_1_346__00555_ (.A(clknet_level_0_1_345__00555_),
    .Z(clknet_level_1_1_346__00555_));
 BUF_X4 clkbuf_level_2_1_347__00555_ (.A(clknet_level_1_1_346__00555_),
    .Z(clknet_level_2_1_347__00555_));
 BUF_X4 clkbuf_level_0_1_448__00555_ (.A(clknet_3_3__leaf__00555_),
    .Z(clknet_level_0_1_448__00555_));
 BUF_X4 clkbuf_level_1_1_449__00555_ (.A(clknet_level_0_1_448__00555_),
    .Z(clknet_level_1_1_449__00555_));
 BUF_X4 clkbuf_level_2_1_450__00555_ (.A(clknet_level_1_1_449__00555_),
    .Z(clknet_level_2_1_450__00555_));
 BUF_X4 clkbuf_level_0_1_551__00555_ (.A(clknet_3_4__leaf__00555_),
    .Z(clknet_level_0_1_551__00555_));
 BUF_X4 clkbuf_level_1_1_552__00555_ (.A(clknet_level_0_1_551__00555_),
    .Z(clknet_level_1_1_552__00555_));
 BUF_X4 clkbuf_level_2_1_553__00555_ (.A(clknet_level_1_1_552__00555_),
    .Z(clknet_level_2_1_553__00555_));
 BUF_X4 clkbuf_level_0_1_654__00555_ (.A(clknet_3_5__leaf__00555_),
    .Z(clknet_level_0_1_654__00555_));
 BUF_X4 clkbuf_level_1_1_655__00555_ (.A(clknet_level_0_1_654__00555_),
    .Z(clknet_level_1_1_655__00555_));
 BUF_X4 clkbuf_level_2_1_656__00555_ (.A(clknet_level_1_1_655__00555_),
    .Z(clknet_level_2_1_656__00555_));
 BUF_X4 clkbuf_level_0_1_757__00555_ (.A(clknet_3_6__leaf__00555_),
    .Z(clknet_level_0_1_757__00555_));
 BUF_X4 clkbuf_level_1_1_758__00555_ (.A(clknet_level_0_1_757__00555_),
    .Z(clknet_level_1_1_758__00555_));
 BUF_X4 clkbuf_level_2_1_759__00555_ (.A(clknet_level_1_1_758__00555_),
    .Z(clknet_level_2_1_759__00555_));
 BUF_X4 clkbuf_level_0_1_860__00555_ (.A(clknet_3_7__leaf__00555_),
    .Z(clknet_level_0_1_860__00555_));
 BUF_X4 clkbuf_level_1_1_861__00555_ (.A(clknet_level_0_1_860__00555_),
    .Z(clknet_level_1_1_861__00555_));
 BUF_X4 clkbuf_level_2_1_862__00555_ (.A(clknet_level_1_1_861__00555_),
    .Z(clknet_level_2_1_862__00555_));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__8.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ));
 BUF_X4 clkbuf_0__00558_ (.A(_00558_),
    .Z(clknet_0__00558_));
 BUF_X4 clkbuf_3_0__f__00558_ (.A(clknet_0__00558_),
    .Z(clknet_3_0__leaf__00558_));
 BUF_X4 clkbuf_3_1__f__00558_ (.A(clknet_0__00558_),
    .Z(clknet_3_1__leaf__00558_));
 BUF_X4 clkbuf_3_2__f__00558_ (.A(clknet_0__00558_),
    .Z(clknet_3_2__leaf__00558_));
 BUF_X4 clkbuf_3_3__f__00558_ (.A(clknet_0__00558_),
    .Z(clknet_3_3__leaf__00558_));
 BUF_X4 clkbuf_3_4__f__00558_ (.A(clknet_0__00558_),
    .Z(clknet_3_4__leaf__00558_));
 BUF_X4 clkbuf_3_5__f__00558_ (.A(clknet_0__00558_),
    .Z(clknet_3_5__leaf__00558_));
 BUF_X4 clkbuf_3_6__f__00558_ (.A(clknet_0__00558_),
    .Z(clknet_3_6__leaf__00558_));
 BUF_X4 clkbuf_3_7__f__00558_ (.A(clknet_0__00558_),
    .Z(clknet_3_7__leaf__00558_));
 BUF_X4 clkbuf_level_0_1_163__00558_ (.A(clknet_3_0__leaf__00558_),
    .Z(clknet_level_0_1_163__00558_));
 BUF_X4 clkbuf_level_1_1_164__00558_ (.A(clknet_level_0_1_163__00558_),
    .Z(clknet_level_1_1_164__00558_));
 BUF_X4 clkbuf_level_2_1_165__00558_ (.A(clknet_level_1_1_164__00558_),
    .Z(clknet_level_2_1_165__00558_));
 BUF_X4 clkbuf_level_0_1_266__00558_ (.A(clknet_3_1__leaf__00558_),
    .Z(clknet_level_0_1_266__00558_));
 BUF_X4 clkbuf_level_1_1_267__00558_ (.A(clknet_level_0_1_266__00558_),
    .Z(clknet_level_1_1_267__00558_));
 BUF_X4 clkbuf_level_2_1_268__00558_ (.A(clknet_level_1_1_267__00558_),
    .Z(clknet_level_2_1_268__00558_));
 BUF_X4 clkbuf_level_0_1_369__00558_ (.A(clknet_3_2__leaf__00558_),
    .Z(clknet_level_0_1_369__00558_));
 BUF_X4 clkbuf_level_1_1_370__00558_ (.A(clknet_level_0_1_369__00558_),
    .Z(clknet_level_1_1_370__00558_));
 BUF_X4 clkbuf_level_2_1_371__00558_ (.A(clknet_level_1_1_370__00558_),
    .Z(clknet_level_2_1_371__00558_));
 BUF_X4 clkbuf_level_0_1_472__00558_ (.A(clknet_3_3__leaf__00558_),
    .Z(clknet_level_0_1_472__00558_));
 BUF_X4 clkbuf_level_1_1_473__00558_ (.A(clknet_level_0_1_472__00558_),
    .Z(clknet_level_1_1_473__00558_));
 BUF_X4 clkbuf_level_2_1_474__00558_ (.A(clknet_level_1_1_473__00558_),
    .Z(clknet_level_2_1_474__00558_));
 BUF_X4 clkbuf_level_0_1_575__00558_ (.A(clknet_3_4__leaf__00558_),
    .Z(clknet_level_0_1_575__00558_));
 BUF_X4 clkbuf_level_1_1_576__00558_ (.A(clknet_level_0_1_575__00558_),
    .Z(clknet_level_1_1_576__00558_));
 BUF_X4 clkbuf_level_2_1_577__00558_ (.A(clknet_level_1_1_576__00558_),
    .Z(clknet_level_2_1_577__00558_));
 BUF_X4 clkbuf_level_0_1_678__00558_ (.A(clknet_3_5__leaf__00558_),
    .Z(clknet_level_0_1_678__00558_));
 BUF_X4 clkbuf_level_1_1_679__00558_ (.A(clknet_level_0_1_678__00558_),
    .Z(clknet_level_1_1_679__00558_));
 BUF_X4 clkbuf_level_2_1_680__00558_ (.A(clknet_level_1_1_679__00558_),
    .Z(clknet_level_2_1_680__00558_));
 BUF_X4 clkbuf_level_0_1_781__00558_ (.A(clknet_3_6__leaf__00558_),
    .Z(clknet_level_0_1_781__00558_));
 BUF_X4 clkbuf_level_1_1_782__00558_ (.A(clknet_level_0_1_781__00558_),
    .Z(clknet_level_1_1_782__00558_));
 BUF_X4 clkbuf_level_2_1_783__00558_ (.A(clknet_level_1_1_782__00558_),
    .Z(clknet_level_2_1_783__00558_));
 BUF_X4 clkbuf_level_0_1_884__00558_ (.A(clknet_3_7__leaf__00558_),
    .Z(clknet_level_0_1_884__00558_));
 BUF_X4 clkbuf_level_1_1_885__00558_ (.A(clknet_level_0_1_884__00558_),
    .Z(clknet_level_1_1_885__00558_));
 BUF_X4 clkbuf_level_2_1_886__00558_ (.A(clknet_level_1_1_885__00558_),
    .Z(clknet_level_2_1_886__00558_));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__7.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ));
 BUF_X4 clkbuf_0__00561_ (.A(_00561_),
    .Z(clknet_0__00561_));
 BUF_X4 clkbuf_3_0__f__00561_ (.A(clknet_0__00561_),
    .Z(clknet_3_0__leaf__00561_));
 BUF_X4 clkbuf_3_1__f__00561_ (.A(clknet_0__00561_),
    .Z(clknet_3_1__leaf__00561_));
 BUF_X4 clkbuf_3_2__f__00561_ (.A(clknet_0__00561_),
    .Z(clknet_3_2__leaf__00561_));
 BUF_X4 clkbuf_3_3__f__00561_ (.A(clknet_0__00561_),
    .Z(clknet_3_3__leaf__00561_));
 BUF_X4 clkbuf_3_4__f__00561_ (.A(clknet_0__00561_),
    .Z(clknet_3_4__leaf__00561_));
 BUF_X4 clkbuf_3_5__f__00561_ (.A(clknet_0__00561_),
    .Z(clknet_3_5__leaf__00561_));
 BUF_X4 clkbuf_3_6__f__00561_ (.A(clknet_0__00561_),
    .Z(clknet_3_6__leaf__00561_));
 BUF_X4 clkbuf_3_7__f__00561_ (.A(clknet_0__00561_),
    .Z(clknet_3_7__leaf__00561_));
 BUF_X4 clkbuf_level_0_1_187__00561_ (.A(clknet_3_0__leaf__00561_),
    .Z(clknet_level_0_1_187__00561_));
 BUF_X4 clkbuf_level_1_1_188__00561_ (.A(clknet_level_0_1_187__00561_),
    .Z(clknet_level_1_1_188__00561_));
 BUF_X4 clkbuf_level_2_1_189__00561_ (.A(clknet_level_1_1_188__00561_),
    .Z(clknet_level_2_1_189__00561_));
 BUF_X4 clkbuf_level_0_1_290__00561_ (.A(clknet_3_1__leaf__00561_),
    .Z(clknet_level_0_1_290__00561_));
 BUF_X4 clkbuf_level_1_1_291__00561_ (.A(clknet_level_0_1_290__00561_),
    .Z(clknet_level_1_1_291__00561_));
 BUF_X4 clkbuf_level_2_1_292__00561_ (.A(clknet_level_1_1_291__00561_),
    .Z(clknet_level_2_1_292__00561_));
 BUF_X4 clkbuf_level_0_1_393__00561_ (.A(clknet_3_2__leaf__00561_),
    .Z(clknet_level_0_1_393__00561_));
 BUF_X4 clkbuf_level_1_1_394__00561_ (.A(clknet_level_0_1_393__00561_),
    .Z(clknet_level_1_1_394__00561_));
 BUF_X4 clkbuf_level_2_1_395__00561_ (.A(clknet_level_1_1_394__00561_),
    .Z(clknet_level_2_1_395__00561_));
 BUF_X4 clkbuf_level_0_1_496__00561_ (.A(clknet_3_3__leaf__00561_),
    .Z(clknet_level_0_1_496__00561_));
 BUF_X4 clkbuf_level_1_1_497__00561_ (.A(clknet_level_0_1_496__00561_),
    .Z(clknet_level_1_1_497__00561_));
 BUF_X4 clkbuf_level_2_1_498__00561_ (.A(clknet_level_1_1_497__00561_),
    .Z(clknet_level_2_1_498__00561_));
 BUF_X4 clkbuf_level_0_1_599__00561_ (.A(clknet_3_4__leaf__00561_),
    .Z(clknet_level_0_1_599__00561_));
 BUF_X4 clkbuf_level_1_1_5100__00561_ (.A(clknet_level_0_1_599__00561_),
    .Z(clknet_level_1_1_5100__00561_));
 BUF_X4 clkbuf_level_2_1_5101__00561_ (.A(clknet_level_1_1_5100__00561_),
    .Z(clknet_level_2_1_5101__00561_));
 BUF_X4 clkbuf_level_0_1_6102__00561_ (.A(clknet_3_5__leaf__00561_),
    .Z(clknet_level_0_1_6102__00561_));
 BUF_X4 clkbuf_level_1_1_6103__00561_ (.A(clknet_level_0_1_6102__00561_),
    .Z(clknet_level_1_1_6103__00561_));
 BUF_X4 clkbuf_level_2_1_6104__00561_ (.A(clknet_level_1_1_6103__00561_),
    .Z(clknet_level_2_1_6104__00561_));
 BUF_X4 clkbuf_level_0_1_7105__00561_ (.A(clknet_3_6__leaf__00561_),
    .Z(clknet_level_0_1_7105__00561_));
 BUF_X4 clkbuf_level_1_1_7106__00561_ (.A(clknet_level_0_1_7105__00561_),
    .Z(clknet_level_1_1_7106__00561_));
 BUF_X4 clkbuf_level_2_1_7107__00561_ (.A(clknet_level_1_1_7106__00561_),
    .Z(clknet_level_2_1_7107__00561_));
 BUF_X4 clkbuf_level_0_1_8108__00561_ (.A(clknet_3_7__leaf__00561_),
    .Z(clknet_level_0_1_8108__00561_));
 BUF_X4 clkbuf_level_1_1_8109__00561_ (.A(clknet_level_0_1_8108__00561_),
    .Z(clknet_level_1_1_8109__00561_));
 BUF_X4 clkbuf_level_2_1_8110__00561_ (.A(clknet_level_1_1_8109__00561_),
    .Z(clknet_level_2_1_8110__00561_));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__6.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ));
 BUF_X4 clkbuf_0__00564_ (.A(_00564_),
    .Z(clknet_0__00564_));
 BUF_X4 clkbuf_3_0__f__00564_ (.A(clknet_0__00564_),
    .Z(clknet_3_0__leaf__00564_));
 BUF_X4 clkbuf_3_1__f__00564_ (.A(clknet_0__00564_),
    .Z(clknet_3_1__leaf__00564_));
 BUF_X4 clkbuf_3_2__f__00564_ (.A(clknet_0__00564_),
    .Z(clknet_3_2__leaf__00564_));
 BUF_X4 clkbuf_3_3__f__00564_ (.A(clknet_0__00564_),
    .Z(clknet_3_3__leaf__00564_));
 BUF_X4 clkbuf_3_4__f__00564_ (.A(clknet_0__00564_),
    .Z(clknet_3_4__leaf__00564_));
 BUF_X4 clkbuf_3_5__f__00564_ (.A(clknet_0__00564_),
    .Z(clknet_3_5__leaf__00564_));
 BUF_X4 clkbuf_3_6__f__00564_ (.A(clknet_0__00564_),
    .Z(clknet_3_6__leaf__00564_));
 BUF_X4 clkbuf_3_7__f__00564_ (.A(clknet_0__00564_),
    .Z(clknet_3_7__leaf__00564_));
 BUF_X4 clkbuf_level_0_1_1243__00564_ (.A(clknet_3_0__leaf__00564_),
    .Z(clknet_level_0_1_1243__00564_));
 BUF_X4 clkbuf_level_1_1_1244__00564_ (.A(clknet_level_0_1_1243__00564_),
    .Z(clknet_level_1_1_1244__00564_));
 BUF_X4 clkbuf_level_2_1_1245__00564_ (.A(clknet_level_1_1_1244__00564_),
    .Z(clknet_level_2_1_1245__00564_));
 BUF_X4 clkbuf_level_0_1_2246__00564_ (.A(clknet_3_1__leaf__00564_),
    .Z(clknet_level_0_1_2246__00564_));
 BUF_X4 clkbuf_level_1_1_2247__00564_ (.A(clknet_level_0_1_2246__00564_),
    .Z(clknet_level_1_1_2247__00564_));
 BUF_X4 clkbuf_level_2_1_2248__00564_ (.A(clknet_level_1_1_2247__00564_),
    .Z(clknet_level_2_1_2248__00564_));
 BUF_X4 clkbuf_level_0_1_3249__00564_ (.A(clknet_3_2__leaf__00564_),
    .Z(clknet_level_0_1_3249__00564_));
 BUF_X4 clkbuf_level_1_1_3250__00564_ (.A(clknet_level_0_1_3249__00564_),
    .Z(clknet_level_1_1_3250__00564_));
 BUF_X4 clkbuf_level_2_1_3251__00564_ (.A(clknet_level_1_1_3250__00564_),
    .Z(clknet_level_2_1_3251__00564_));
 BUF_X4 clkbuf_level_0_1_4252__00564_ (.A(clknet_3_3__leaf__00564_),
    .Z(clknet_level_0_1_4252__00564_));
 BUF_X4 clkbuf_level_1_1_4253__00564_ (.A(clknet_level_0_1_4252__00564_),
    .Z(clknet_level_1_1_4253__00564_));
 BUF_X4 clkbuf_level_2_1_4254__00564_ (.A(clknet_level_1_1_4253__00564_),
    .Z(clknet_level_2_1_4254__00564_));
 BUF_X4 clkbuf_level_0_1_5255__00564_ (.A(clknet_3_4__leaf__00564_),
    .Z(clknet_level_0_1_5255__00564_));
 BUF_X4 clkbuf_level_1_1_5256__00564_ (.A(clknet_level_0_1_5255__00564_),
    .Z(clknet_level_1_1_5256__00564_));
 BUF_X4 clkbuf_level_2_1_5257__00564_ (.A(clknet_level_1_1_5256__00564_),
    .Z(clknet_level_2_1_5257__00564_));
 BUF_X4 clkbuf_level_0_1_6258__00564_ (.A(clknet_3_5__leaf__00564_),
    .Z(clknet_level_0_1_6258__00564_));
 BUF_X4 clkbuf_level_1_1_6259__00564_ (.A(clknet_level_0_1_6258__00564_),
    .Z(clknet_level_1_1_6259__00564_));
 BUF_X4 clkbuf_level_2_1_6260__00564_ (.A(clknet_level_1_1_6259__00564_),
    .Z(clknet_level_2_1_6260__00564_));
 BUF_X4 clkbuf_level_0_1_7261__00564_ (.A(clknet_3_6__leaf__00564_),
    .Z(clknet_level_0_1_7261__00564_));
 BUF_X4 clkbuf_level_1_1_7262__00564_ (.A(clknet_level_0_1_7261__00564_),
    .Z(clknet_level_1_1_7262__00564_));
 BUF_X4 clkbuf_level_2_1_7263__00564_ (.A(clknet_level_1_1_7262__00564_),
    .Z(clknet_level_2_1_7263__00564_));
 BUF_X4 clkbuf_level_0_1_8264__00564_ (.A(clknet_3_7__leaf__00564_),
    .Z(clknet_level_0_1_8264__00564_));
 BUF_X4 clkbuf_level_1_1_8265__00564_ (.A(clknet_level_0_1_8264__00564_),
    .Z(clknet_level_1_1_8265__00564_));
 BUF_X4 clkbuf_level_2_1_8266__00564_ (.A(clknet_level_1_1_8265__00564_),
    .Z(clknet_level_2_1_8266__00564_));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__5.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ));
 BUF_X4 clkbuf_0__00567_ (.A(_00567_),
    .Z(clknet_0__00567_));
 BUF_X4 clkbuf_3_0__f__00567_ (.A(clknet_0__00567_),
    .Z(clknet_3_0__leaf__00567_));
 BUF_X4 clkbuf_3_1__f__00567_ (.A(clknet_0__00567_),
    .Z(clknet_3_1__leaf__00567_));
 BUF_X4 clkbuf_3_2__f__00567_ (.A(clknet_0__00567_),
    .Z(clknet_3_2__leaf__00567_));
 BUF_X4 clkbuf_3_3__f__00567_ (.A(clknet_0__00567_),
    .Z(clknet_3_3__leaf__00567_));
 BUF_X4 clkbuf_3_4__f__00567_ (.A(clknet_0__00567_),
    .Z(clknet_3_4__leaf__00567_));
 BUF_X4 clkbuf_3_5__f__00567_ (.A(clknet_0__00567_),
    .Z(clknet_3_5__leaf__00567_));
 BUF_X4 clkbuf_3_6__f__00567_ (.A(clknet_0__00567_),
    .Z(clknet_3_6__leaf__00567_));
 BUF_X4 clkbuf_3_7__f__00567_ (.A(clknet_0__00567_),
    .Z(clknet_3_7__leaf__00567_));
 BUF_X4 clkbuf_level_0_1_1189__00567_ (.A(clknet_3_0__leaf__00567_),
    .Z(clknet_level_0_1_1189__00567_));
 BUF_X4 clkbuf_level_1_1_1190__00567_ (.A(clknet_level_0_1_1189__00567_),
    .Z(clknet_level_1_1_1190__00567_));
 BUF_X4 clkbuf_level_2_1_1191__00567_ (.A(clknet_level_1_1_1190__00567_),
    .Z(clknet_level_2_1_1191__00567_));
 BUF_X4 clkbuf_level_0_1_2192__00567_ (.A(clknet_3_1__leaf__00567_),
    .Z(clknet_level_0_1_2192__00567_));
 BUF_X4 clkbuf_level_1_1_2193__00567_ (.A(clknet_level_0_1_2192__00567_),
    .Z(clknet_level_1_1_2193__00567_));
 BUF_X4 clkbuf_level_2_1_2194__00567_ (.A(clknet_level_1_1_2193__00567_),
    .Z(clknet_level_2_1_2194__00567_));
 BUF_X4 clkbuf_level_0_1_3195__00567_ (.A(clknet_3_2__leaf__00567_),
    .Z(clknet_level_0_1_3195__00567_));
 BUF_X4 clkbuf_level_1_1_3196__00567_ (.A(clknet_level_0_1_3195__00567_),
    .Z(clknet_level_1_1_3196__00567_));
 BUF_X4 clkbuf_level_2_1_3197__00567_ (.A(clknet_level_1_1_3196__00567_),
    .Z(clknet_level_2_1_3197__00567_));
 BUF_X4 clkbuf_level_0_1_4198__00567_ (.A(clknet_3_3__leaf__00567_),
    .Z(clknet_level_0_1_4198__00567_));
 BUF_X4 clkbuf_level_1_1_4199__00567_ (.A(clknet_level_0_1_4198__00567_),
    .Z(clknet_level_1_1_4199__00567_));
 BUF_X4 clkbuf_level_2_1_4200__00567_ (.A(clknet_level_1_1_4199__00567_),
    .Z(clknet_level_2_1_4200__00567_));
 BUF_X4 clkbuf_level_0_1_5201__00567_ (.A(clknet_3_4__leaf__00567_),
    .Z(clknet_level_0_1_5201__00567_));
 BUF_X4 clkbuf_level_1_1_5202__00567_ (.A(clknet_level_0_1_5201__00567_),
    .Z(clknet_level_1_1_5202__00567_));
 BUF_X4 clkbuf_level_2_1_5203__00567_ (.A(clknet_level_1_1_5202__00567_),
    .Z(clknet_level_2_1_5203__00567_));
 BUF_X4 clkbuf_level_0_1_6204__00567_ (.A(clknet_3_5__leaf__00567_),
    .Z(clknet_level_0_1_6204__00567_));
 BUF_X4 clkbuf_level_1_1_6205__00567_ (.A(clknet_level_0_1_6204__00567_),
    .Z(clknet_level_1_1_6205__00567_));
 BUF_X4 clkbuf_level_2_1_6206__00567_ (.A(clknet_level_1_1_6205__00567_),
    .Z(clknet_level_2_1_6206__00567_));
 BUF_X4 clkbuf_level_0_1_7207__00567_ (.A(clknet_3_6__leaf__00567_),
    .Z(clknet_level_0_1_7207__00567_));
 BUF_X4 clkbuf_level_1_1_7208__00567_ (.A(clknet_level_0_1_7207__00567_),
    .Z(clknet_level_1_1_7208__00567_));
 BUF_X4 clkbuf_level_2_1_7209__00567_ (.A(clknet_level_1_1_7208__00567_),
    .Z(clknet_level_2_1_7209__00567_));
 BUF_X4 clkbuf_level_0_1_8210__00567_ (.A(clknet_3_7__leaf__00567_),
    .Z(clknet_level_0_1_8210__00567_));
 BUF_X4 clkbuf_level_1_1_8211__00567_ (.A(clknet_level_0_1_8210__00567_),
    .Z(clknet_level_1_1_8211__00567_));
 BUF_X4 clkbuf_level_2_1_8212__00567_ (.A(clknet_level_1_1_8211__00567_),
    .Z(clknet_level_2_1_8212__00567_));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__4.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ));
 BUF_X4 clkbuf_0__00570_ (.A(_00570_),
    .Z(clknet_0__00570_));
 BUF_X4 clkbuf_3_0__f__00570_ (.A(clknet_0__00570_),
    .Z(clknet_3_0__leaf__00570_));
 BUF_X4 clkbuf_3_1__f__00570_ (.A(clknet_0__00570_),
    .Z(clknet_3_1__leaf__00570_));
 BUF_X4 clkbuf_3_2__f__00570_ (.A(clknet_0__00570_),
    .Z(clknet_3_2__leaf__00570_));
 BUF_X4 clkbuf_3_3__f__00570_ (.A(clknet_0__00570_),
    .Z(clknet_3_3__leaf__00570_));
 BUF_X4 clkbuf_3_4__f__00570_ (.A(clknet_0__00570_),
    .Z(clknet_3_4__leaf__00570_));
 BUF_X4 clkbuf_3_5__f__00570_ (.A(clknet_0__00570_),
    .Z(clknet_3_5__leaf__00570_));
 BUF_X4 clkbuf_3_6__f__00570_ (.A(clknet_0__00570_),
    .Z(clknet_3_6__leaf__00570_));
 BUF_X4 clkbuf_3_7__f__00570_ (.A(clknet_0__00570_),
    .Z(clknet_3_7__leaf__00570_));
 BUF_X4 clkbuf_level_0_1_1267__00570_ (.A(clknet_3_0__leaf__00570_),
    .Z(clknet_level_0_1_1267__00570_));
 BUF_X4 clkbuf_level_1_1_1268__00570_ (.A(clknet_level_0_1_1267__00570_),
    .Z(clknet_level_1_1_1268__00570_));
 BUF_X4 clkbuf_level_2_1_1269__00570_ (.A(clknet_level_1_1_1268__00570_),
    .Z(clknet_level_2_1_1269__00570_));
 BUF_X4 clkbuf_level_0_1_2270__00570_ (.A(clknet_3_1__leaf__00570_),
    .Z(clknet_level_0_1_2270__00570_));
 BUF_X4 clkbuf_level_1_1_2271__00570_ (.A(clknet_level_0_1_2270__00570_),
    .Z(clknet_level_1_1_2271__00570_));
 BUF_X4 clkbuf_level_2_1_2272__00570_ (.A(clknet_level_1_1_2271__00570_),
    .Z(clknet_level_2_1_2272__00570_));
 BUF_X4 clkbuf_level_0_1_3273__00570_ (.A(clknet_3_2__leaf__00570_),
    .Z(clknet_level_0_1_3273__00570_));
 BUF_X4 clkbuf_level_1_1_3274__00570_ (.A(clknet_level_0_1_3273__00570_),
    .Z(clknet_level_1_1_3274__00570_));
 BUF_X4 clkbuf_level_2_1_3275__00570_ (.A(clknet_level_1_1_3274__00570_),
    .Z(clknet_level_2_1_3275__00570_));
 BUF_X4 clkbuf_level_0_1_4276__00570_ (.A(clknet_3_3__leaf__00570_),
    .Z(clknet_level_0_1_4276__00570_));
 BUF_X4 clkbuf_level_1_1_4277__00570_ (.A(clknet_level_0_1_4276__00570_),
    .Z(clknet_level_1_1_4277__00570_));
 BUF_X4 clkbuf_level_2_1_4278__00570_ (.A(clknet_level_1_1_4277__00570_),
    .Z(clknet_level_2_1_4278__00570_));
 BUF_X4 clkbuf_level_0_1_5279__00570_ (.A(clknet_3_4__leaf__00570_),
    .Z(clknet_level_0_1_5279__00570_));
 BUF_X4 clkbuf_level_1_1_5280__00570_ (.A(clknet_level_0_1_5279__00570_),
    .Z(clknet_level_1_1_5280__00570_));
 BUF_X4 clkbuf_level_2_1_5281__00570_ (.A(clknet_level_1_1_5280__00570_),
    .Z(clknet_level_2_1_5281__00570_));
 BUF_X4 clkbuf_level_0_1_6282__00570_ (.A(clknet_3_5__leaf__00570_),
    .Z(clknet_level_0_1_6282__00570_));
 BUF_X4 clkbuf_level_1_1_6283__00570_ (.A(clknet_level_0_1_6282__00570_),
    .Z(clknet_level_1_1_6283__00570_));
 BUF_X4 clkbuf_level_2_1_6284__00570_ (.A(clknet_level_1_1_6283__00570_),
    .Z(clknet_level_2_1_6284__00570_));
 BUF_X4 clkbuf_level_0_1_7285__00570_ (.A(clknet_3_6__leaf__00570_),
    .Z(clknet_level_0_1_7285__00570_));
 BUF_X4 clkbuf_level_1_1_7286__00570_ (.A(clknet_level_0_1_7285__00570_),
    .Z(clknet_level_1_1_7286__00570_));
 BUF_X4 clkbuf_level_2_1_7287__00570_ (.A(clknet_level_1_1_7286__00570_),
    .Z(clknet_level_2_1_7287__00570_));
 BUF_X4 clkbuf_level_0_1_8288__00570_ (.A(clknet_3_7__leaf__00570_),
    .Z(clknet_level_0_1_8288__00570_));
 BUF_X4 clkbuf_level_1_1_8289__00570_ (.A(clknet_level_0_1_8288__00570_),
    .Z(clknet_level_1_1_8289__00570_));
 BUF_X4 clkbuf_level_2_1_8290__00570_ (.A(clknet_level_1_1_8289__00570_),
    .Z(clknet_level_2_1_8290__00570_));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__3.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ));
 BUF_X4 clkbuf_0__00573_ (.A(_00573_),
    .Z(clknet_0__00573_));
 BUF_X4 clkbuf_3_0__f__00573_ (.A(clknet_0__00573_),
    .Z(clknet_3_0__leaf__00573_));
 BUF_X4 clkbuf_3_1__f__00573_ (.A(clknet_0__00573_),
    .Z(clknet_3_1__leaf__00573_));
 BUF_X4 clkbuf_3_2__f__00573_ (.A(clknet_0__00573_),
    .Z(clknet_3_2__leaf__00573_));
 BUF_X4 clkbuf_3_3__f__00573_ (.A(clknet_0__00573_),
    .Z(clknet_3_3__leaf__00573_));
 BUF_X4 clkbuf_3_4__f__00573_ (.A(clknet_0__00573_),
    .Z(clknet_3_4__leaf__00573_));
 BUF_X4 clkbuf_3_5__f__00573_ (.A(clknet_0__00573_),
    .Z(clknet_3_5__leaf__00573_));
 BUF_X4 clkbuf_3_6__f__00573_ (.A(clknet_0__00573_),
    .Z(clknet_3_6__leaf__00573_));
 BUF_X4 clkbuf_3_7__f__00573_ (.A(clknet_0__00573_),
    .Z(clknet_3_7__leaf__00573_));
 BUF_X4 clkbuf_level_0_1_1291__00573_ (.A(clknet_3_0__leaf__00573_),
    .Z(clknet_level_0_1_1291__00573_));
 BUF_X4 clkbuf_level_1_1_1292__00573_ (.A(clknet_level_0_1_1291__00573_),
    .Z(clknet_level_1_1_1292__00573_));
 BUF_X4 clkbuf_level_2_1_1293__00573_ (.A(clknet_level_1_1_1292__00573_),
    .Z(clknet_level_2_1_1293__00573_));
 BUF_X4 clkbuf_level_0_1_2294__00573_ (.A(clknet_3_1__leaf__00573_),
    .Z(clknet_level_0_1_2294__00573_));
 BUF_X4 clkbuf_level_1_1_2295__00573_ (.A(clknet_level_0_1_2294__00573_),
    .Z(clknet_level_1_1_2295__00573_));
 BUF_X4 clkbuf_level_2_1_2296__00573_ (.A(clknet_level_1_1_2295__00573_),
    .Z(clknet_level_2_1_2296__00573_));
 BUF_X4 clkbuf_level_0_1_3297__00573_ (.A(clknet_3_2__leaf__00573_),
    .Z(clknet_level_0_1_3297__00573_));
 BUF_X4 clkbuf_level_1_1_3298__00573_ (.A(clknet_level_0_1_3297__00573_),
    .Z(clknet_level_1_1_3298__00573_));
 BUF_X4 clkbuf_level_2_1_3299__00573_ (.A(clknet_level_1_1_3298__00573_),
    .Z(clknet_level_2_1_3299__00573_));
 BUF_X4 clkbuf_level_0_1_4300__00573_ (.A(clknet_3_3__leaf__00573_),
    .Z(clknet_level_0_1_4300__00573_));
 BUF_X4 clkbuf_level_1_1_4301__00573_ (.A(clknet_level_0_1_4300__00573_),
    .Z(clknet_level_1_1_4301__00573_));
 BUF_X4 clkbuf_level_2_1_4302__00573_ (.A(clknet_level_1_1_4301__00573_),
    .Z(clknet_level_2_1_4302__00573_));
 BUF_X4 clkbuf_level_0_1_5303__00573_ (.A(clknet_3_4__leaf__00573_),
    .Z(clknet_level_0_1_5303__00573_));
 BUF_X4 clkbuf_level_1_1_5304__00573_ (.A(clknet_level_0_1_5303__00573_),
    .Z(clknet_level_1_1_5304__00573_));
 BUF_X4 clkbuf_level_2_1_5305__00573_ (.A(clknet_level_1_1_5304__00573_),
    .Z(clknet_level_2_1_5305__00573_));
 BUF_X4 clkbuf_level_0_1_6306__00573_ (.A(clknet_3_5__leaf__00573_),
    .Z(clknet_level_0_1_6306__00573_));
 BUF_X4 clkbuf_level_1_1_6307__00573_ (.A(clknet_level_0_1_6306__00573_),
    .Z(clknet_level_1_1_6307__00573_));
 BUF_X4 clkbuf_level_2_1_6308__00573_ (.A(clknet_level_1_1_6307__00573_),
    .Z(clknet_level_2_1_6308__00573_));
 BUF_X4 clkbuf_level_0_1_7309__00573_ (.A(clknet_3_6__leaf__00573_),
    .Z(clknet_level_0_1_7309__00573_));
 BUF_X4 clkbuf_level_1_1_7310__00573_ (.A(clknet_level_0_1_7309__00573_),
    .Z(clknet_level_1_1_7310__00573_));
 BUF_X4 clkbuf_level_2_1_7311__00573_ (.A(clknet_level_1_1_7310__00573_),
    .Z(clknet_level_2_1_7311__00573_));
 BUF_X4 clkbuf_level_0_1_8312__00573_ (.A(clknet_3_7__leaf__00573_),
    .Z(clknet_level_0_1_8312__00573_));
 BUF_X4 clkbuf_level_1_1_8313__00573_ (.A(clknet_level_0_1_8312__00573_),
    .Z(clknet_level_1_1_8313__00573_));
 BUF_X4 clkbuf_level_2_1_8314__00573_ (.A(clknet_level_1_1_8313__00573_),
    .Z(clknet_level_2_1_8314__00573_));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__2.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ));
 BUF_X4 clkbuf_0__00576_ (.A(_00576_),
    .Z(clknet_0__00576_));
 BUF_X4 clkbuf_3_0__f__00576_ (.A(clknet_0__00576_),
    .Z(clknet_3_0__leaf__00576_));
 BUF_X4 clkbuf_3_1__f__00576_ (.A(clknet_0__00576_),
    .Z(clknet_3_1__leaf__00576_));
 BUF_X4 clkbuf_3_2__f__00576_ (.A(clknet_0__00576_),
    .Z(clknet_3_2__leaf__00576_));
 BUF_X4 clkbuf_3_3__f__00576_ (.A(clknet_0__00576_),
    .Z(clknet_3_3__leaf__00576_));
 BUF_X4 clkbuf_3_4__f__00576_ (.A(clknet_0__00576_),
    .Z(clknet_3_4__leaf__00576_));
 BUF_X4 clkbuf_3_5__f__00576_ (.A(clknet_0__00576_),
    .Z(clknet_3_5__leaf__00576_));
 BUF_X4 clkbuf_3_6__f__00576_ (.A(clknet_0__00576_),
    .Z(clknet_3_6__leaf__00576_));
 BUF_X4 clkbuf_3_7__f__00576_ (.A(clknet_0__00576_),
    .Z(clknet_3_7__leaf__00576_));
 BUF_X4 clkbuf_level_0_1_1369__00576_ (.A(clknet_3_0__leaf__00576_),
    .Z(clknet_level_0_1_1369__00576_));
 BUF_X4 clkbuf_level_1_1_1370__00576_ (.A(clknet_level_0_1_1369__00576_),
    .Z(clknet_level_1_1_1370__00576_));
 BUF_X4 clkbuf_level_2_1_1371__00576_ (.A(clknet_level_1_1_1370__00576_),
    .Z(clknet_level_2_1_1371__00576_));
 BUF_X4 clkbuf_level_0_1_2372__00576_ (.A(clknet_3_1__leaf__00576_),
    .Z(clknet_level_0_1_2372__00576_));
 BUF_X4 clkbuf_level_1_1_2373__00576_ (.A(clknet_level_0_1_2372__00576_),
    .Z(clknet_level_1_1_2373__00576_));
 BUF_X4 clkbuf_level_2_1_2374__00576_ (.A(clknet_level_1_1_2373__00576_),
    .Z(clknet_level_2_1_2374__00576_));
 BUF_X4 clkbuf_level_0_1_3375__00576_ (.A(clknet_3_2__leaf__00576_),
    .Z(clknet_level_0_1_3375__00576_));
 BUF_X4 clkbuf_level_1_1_3376__00576_ (.A(clknet_level_0_1_3375__00576_),
    .Z(clknet_level_1_1_3376__00576_));
 BUF_X4 clkbuf_level_2_1_3377__00576_ (.A(clknet_level_1_1_3376__00576_),
    .Z(clknet_level_2_1_3377__00576_));
 BUF_X4 clkbuf_level_0_1_4378__00576_ (.A(clknet_3_3__leaf__00576_),
    .Z(clknet_level_0_1_4378__00576_));
 BUF_X4 clkbuf_level_1_1_4379__00576_ (.A(clknet_level_0_1_4378__00576_),
    .Z(clknet_level_1_1_4379__00576_));
 BUF_X4 clkbuf_level_2_1_4380__00576_ (.A(clknet_level_1_1_4379__00576_),
    .Z(clknet_level_2_1_4380__00576_));
 BUF_X4 clkbuf_level_0_1_5381__00576_ (.A(clknet_3_4__leaf__00576_),
    .Z(clknet_level_0_1_5381__00576_));
 BUF_X4 clkbuf_level_1_1_5382__00576_ (.A(clknet_level_0_1_5381__00576_),
    .Z(clknet_level_1_1_5382__00576_));
 BUF_X4 clkbuf_level_2_1_5383__00576_ (.A(clknet_level_1_1_5382__00576_),
    .Z(clknet_level_2_1_5383__00576_));
 BUF_X4 clkbuf_level_0_1_6384__00576_ (.A(clknet_3_5__leaf__00576_),
    .Z(clknet_level_0_1_6384__00576_));
 BUF_X4 clkbuf_level_1_1_6385__00576_ (.A(clknet_level_0_1_6384__00576_),
    .Z(clknet_level_1_1_6385__00576_));
 BUF_X4 clkbuf_level_2_1_6386__00576_ (.A(clknet_level_1_1_6385__00576_),
    .Z(clknet_level_2_1_6386__00576_));
 BUF_X4 clkbuf_level_0_1_7387__00576_ (.A(clknet_3_6__leaf__00576_),
    .Z(clknet_level_0_1_7387__00576_));
 BUF_X4 clkbuf_level_1_1_7388__00576_ (.A(clknet_level_0_1_7387__00576_),
    .Z(clknet_level_1_1_7388__00576_));
 BUF_X4 clkbuf_level_2_1_7389__00576_ (.A(clknet_level_1_1_7388__00576_),
    .Z(clknet_level_2_1_7389__00576_));
 BUF_X4 clkbuf_level_0_1_8390__00576_ (.A(clknet_3_7__leaf__00576_),
    .Z(clknet_level_0_1_8390__00576_));
 BUF_X4 clkbuf_level_1_1_8391__00576_ (.A(clknet_level_0_1_8390__00576_),
    .Z(clknet_level_1_1_8391__00576_));
 BUF_X4 clkbuf_level_2_1_8392__00576_ (.A(clknet_level_1_1_8391__00576_),
    .Z(clknet_level_2_1_8392__00576_));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__1.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ));
 BUF_X4 clkbuf_0__00579_ (.A(_00579_),
    .Z(clknet_0__00579_));
 BUF_X4 clkbuf_3_0__f__00579_ (.A(clknet_0__00579_),
    .Z(clknet_3_0__leaf__00579_));
 BUF_X4 clkbuf_3_1__f__00579_ (.A(clknet_0__00579_),
    .Z(clknet_3_1__leaf__00579_));
 BUF_X4 clkbuf_3_2__f__00579_ (.A(clknet_0__00579_),
    .Z(clknet_3_2__leaf__00579_));
 BUF_X4 clkbuf_3_3__f__00579_ (.A(clknet_0__00579_),
    .Z(clknet_3_3__leaf__00579_));
 BUF_X4 clkbuf_3_4__f__00579_ (.A(clknet_0__00579_),
    .Z(clknet_3_4__leaf__00579_));
 BUF_X4 clkbuf_3_5__f__00579_ (.A(clknet_0__00579_),
    .Z(clknet_3_5__leaf__00579_));
 BUF_X4 clkbuf_3_6__f__00579_ (.A(clknet_0__00579_),
    .Z(clknet_3_6__leaf__00579_));
 BUF_X4 clkbuf_3_7__f__00579_ (.A(clknet_0__00579_),
    .Z(clknet_3_7__leaf__00579_));
 BUF_X4 clkbuf_level_0_1_1393__00579_ (.A(clknet_3_0__leaf__00579_),
    .Z(clknet_level_0_1_1393__00579_));
 BUF_X4 clkbuf_level_1_1_1394__00579_ (.A(clknet_level_0_1_1393__00579_),
    .Z(clknet_level_1_1_1394__00579_));
 BUF_X4 clkbuf_level_2_1_1395__00579_ (.A(clknet_level_1_1_1394__00579_),
    .Z(clknet_level_2_1_1395__00579_));
 BUF_X4 clkbuf_level_0_1_2396__00579_ (.A(clknet_3_1__leaf__00579_),
    .Z(clknet_level_0_1_2396__00579_));
 BUF_X4 clkbuf_level_1_1_2397__00579_ (.A(clknet_level_0_1_2396__00579_),
    .Z(clknet_level_1_1_2397__00579_));
 BUF_X4 clkbuf_level_2_1_2398__00579_ (.A(clknet_level_1_1_2397__00579_),
    .Z(clknet_level_2_1_2398__00579_));
 BUF_X4 clkbuf_level_0_1_3399__00579_ (.A(clknet_3_2__leaf__00579_),
    .Z(clknet_level_0_1_3399__00579_));
 BUF_X4 clkbuf_level_1_1_3400__00579_ (.A(clknet_level_0_1_3399__00579_),
    .Z(clknet_level_1_1_3400__00579_));
 BUF_X4 clkbuf_level_2_1_3401__00579_ (.A(clknet_level_1_1_3400__00579_),
    .Z(clknet_level_2_1_3401__00579_));
 BUF_X4 clkbuf_level_0_1_4402__00579_ (.A(clknet_3_3__leaf__00579_),
    .Z(clknet_level_0_1_4402__00579_));
 BUF_X4 clkbuf_level_1_1_4403__00579_ (.A(clknet_level_0_1_4402__00579_),
    .Z(clknet_level_1_1_4403__00579_));
 BUF_X4 clkbuf_level_2_1_4404__00579_ (.A(clknet_level_1_1_4403__00579_),
    .Z(clknet_level_2_1_4404__00579_));
 BUF_X4 clkbuf_level_0_1_5405__00579_ (.A(clknet_3_4__leaf__00579_),
    .Z(clknet_level_0_1_5405__00579_));
 BUF_X4 clkbuf_level_1_1_5406__00579_ (.A(clknet_level_0_1_5405__00579_),
    .Z(clknet_level_1_1_5406__00579_));
 BUF_X4 clkbuf_level_2_1_5407__00579_ (.A(clknet_level_1_1_5406__00579_),
    .Z(clknet_level_2_1_5407__00579_));
 BUF_X4 clkbuf_level_0_1_6408__00579_ (.A(clknet_3_5__leaf__00579_),
    .Z(clknet_level_0_1_6408__00579_));
 BUF_X4 clkbuf_level_1_1_6409__00579_ (.A(clknet_level_0_1_6408__00579_),
    .Z(clknet_level_1_1_6409__00579_));
 BUF_X4 clkbuf_level_2_1_6410__00579_ (.A(clknet_level_1_1_6409__00579_),
    .Z(clknet_level_2_1_6410__00579_));
 BUF_X4 clkbuf_level_0_1_7411__00579_ (.A(clknet_3_6__leaf__00579_),
    .Z(clknet_level_0_1_7411__00579_));
 BUF_X4 clkbuf_level_1_1_7412__00579_ (.A(clknet_level_0_1_7411__00579_),
    .Z(clknet_level_1_1_7412__00579_));
 BUF_X4 clkbuf_level_2_1_7413__00579_ (.A(clknet_level_1_1_7412__00579_),
    .Z(clknet_level_2_1_7413__00579_));
 BUF_X4 clkbuf_level_0_1_8414__00579_ (.A(clknet_3_7__leaf__00579_),
    .Z(clknet_level_0_1_8414__00579_));
 BUF_X4 clkbuf_level_1_1_8415__00579_ (.A(clknet_level_0_1_8414__00579_),
    .Z(clknet_level_1_1_8415__00579_));
 BUF_X4 clkbuf_level_2_1_8416__00579_ (.A(clknet_level_1_1_8415__00579_),
    .Z(clknet_level_2_1_8416__00579_));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__19.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__20.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__21.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__22.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__23.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__24.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__25.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__26.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__27.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__28.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__9.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__10.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__11.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__12.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__13.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__14.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__15.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__16.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__17.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__18.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__0.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__1.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__2.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__3.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__4.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__5.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__6.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__7.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__8.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__31.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__30.cg_i.clk_o ));
 BUF_X4 \clkbuf_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o  (.A(\lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Z(\clknet_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_0__f_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Z(\clknet_1_0__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ));
 BUF_X4 \clkbuf_1_1__f_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o  (.A(\clknet_0_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ),
    .Z(\clknet_1_1__leaf_lut.gen_sub_units_scm.__0.sub_unit_i.gen_cg_word_iter.__29.cg_i.clk_o ));
 FILLCELL_X32 FILLER_0_0_1 ();
 FILLCELL_X32 FILLER_0_0_33 ();
 FILLCELL_X32 FILLER_0_0_65 ();
 FILLCELL_X32 FILLER_0_0_97 ();
 FILLCELL_X32 FILLER_0_0_129 ();
 FILLCELL_X32 FILLER_0_0_161 ();
 FILLCELL_X32 FILLER_0_0_193 ();
 FILLCELL_X32 FILLER_0_0_225 ();
 FILLCELL_X32 FILLER_0_0_257 ();
 FILLCELL_X16 FILLER_0_0_289 ();
 FILLCELL_X4 FILLER_0_0_305 ();
 FILLCELL_X2 FILLER_0_0_309 ();
 FILLCELL_X1 FILLER_0_0_311 ();
 FILLCELL_X32 FILLER_0_0_321 ();
 FILLCELL_X16 FILLER_0_0_353 ();
 FILLCELL_X4 FILLER_0_0_369 ();
 FILLCELL_X2 FILLER_0_0_373 ();
 FILLCELL_X1 FILLER_0_0_375 ();
 FILLCELL_X2 FILLER_0_0_425 ();
 FILLCELL_X1 FILLER_0_0_427 ();
 FILLCELL_X2 FILLER_0_0_453 ();
 FILLCELL_X1 FILLER_0_0_455 ();
 FILLCELL_X4 FILLER_0_0_476 ();
 FILLCELL_X4 FILLER_0_0_495 ();
 FILLCELL_X8 FILLER_0_0_508 ();
 FILLCELL_X1 FILLER_0_0_516 ();
 FILLCELL_X2 FILLER_0_0_539 ();
 FILLCELL_X1 FILLER_0_0_541 ();
 FILLCELL_X16 FILLER_0_0_549 ();
 FILLCELL_X8 FILLER_0_0_565 ();
 FILLCELL_X2 FILLER_0_0_573 ();
 FILLCELL_X32 FILLER_0_0_585 ();
 FILLCELL_X4 FILLER_0_0_617 ();
 FILLCELL_X16 FILLER_0_0_632 ();
 FILLCELL_X4 FILLER_0_0_648 ();
 FILLCELL_X1 FILLER_0_0_657 ();
 FILLCELL_X32 FILLER_0_0_663 ();
 FILLCELL_X4 FILLER_0_0_695 ();
 FILLCELL_X2 FILLER_0_0_699 ();
 FILLCELL_X2 FILLER_0_0_716 ();
 FILLCELL_X1 FILLER_0_0_718 ();
 FILLCELL_X2 FILLER_0_0_724 ();
 FILLCELL_X2 FILLER_0_0_748 ();
 FILLCELL_X1 FILLER_0_0_750 ();
 FILLCELL_X32 FILLER_0_0_756 ();
 FILLCELL_X32 FILLER_0_0_788 ();
 FILLCELL_X4 FILLER_0_0_820 ();
 FILLCELL_X1 FILLER_0_0_824 ();
 FILLCELL_X8 FILLER_0_0_855 ();
 FILLCELL_X2 FILLER_0_0_863 ();
 FILLCELL_X8 FILLER_0_0_885 ();
 FILLCELL_X1 FILLER_0_0_893 ();
 FILLCELL_X8 FILLER_0_0_899 ();
 FILLCELL_X4 FILLER_0_0_907 ();
 FILLCELL_X2 FILLER_0_0_911 ();
 FILLCELL_X1 FILLER_0_0_913 ();
 FILLCELL_X4 FILLER_0_0_919 ();
 FILLCELL_X2 FILLER_0_0_923 ();
 FILLCELL_X1 FILLER_0_0_925 ();
 FILLCELL_X4 FILLER_0_0_936 ();
 FILLCELL_X2 FILLER_0_0_957 ();
 FILLCELL_X1 FILLER_0_0_959 ();
 FILLCELL_X4 FILLER_0_0_975 ();
 FILLCELL_X32 FILLER_0_0_994 ();
 FILLCELL_X32 FILLER_0_0_1026 ();
 FILLCELL_X32 FILLER_0_0_1058 ();
 FILLCELL_X32 FILLER_0_0_1090 ();
 FILLCELL_X16 FILLER_0_0_1122 ();
 FILLCELL_X8 FILLER_0_0_1138 ();
 FILLCELL_X2 FILLER_0_0_1146 ();
 FILLCELL_X32 FILLER_0_1_1 ();
 FILLCELL_X32 FILLER_0_1_33 ();
 FILLCELL_X32 FILLER_0_1_65 ();
 FILLCELL_X32 FILLER_0_1_97 ();
 FILLCELL_X32 FILLER_0_1_129 ();
 FILLCELL_X32 FILLER_0_1_161 ();
 FILLCELL_X32 FILLER_0_1_193 ();
 FILLCELL_X32 FILLER_0_1_225 ();
 FILLCELL_X16 FILLER_0_1_257 ();
 FILLCELL_X2 FILLER_0_1_273 ();
 FILLCELL_X4 FILLER_0_1_280 ();
 FILLCELL_X8 FILLER_0_1_291 ();
 FILLCELL_X1 FILLER_0_1_299 ();
 FILLCELL_X8 FILLER_0_1_330 ();
 FILLCELL_X2 FILLER_0_1_348 ();
 FILLCELL_X16 FILLER_0_1_360 ();
 FILLCELL_X8 FILLER_0_1_376 ();
 FILLCELL_X2 FILLER_0_1_384 ();
 FILLCELL_X4 FILLER_0_1_436 ();
 FILLCELL_X1 FILLER_0_1_474 ();
 FILLCELL_X2 FILLER_0_1_509 ();
 FILLCELL_X2 FILLER_0_1_526 ();
 FILLCELL_X1 FILLER_0_1_553 ();
 FILLCELL_X2 FILLER_0_1_569 ();
 FILLCELL_X16 FILLER_0_1_590 ();
 FILLCELL_X4 FILLER_0_1_606 ();
 FILLCELL_X1 FILLER_0_1_620 ();
 FILLCELL_X1 FILLER_0_1_630 ();
 FILLCELL_X2 FILLER_0_1_674 ();
 FILLCELL_X2 FILLER_0_1_696 ();
 FILLCELL_X1 FILLER_0_1_698 ();
 FILLCELL_X4 FILLER_0_1_704 ();
 FILLCELL_X2 FILLER_0_1_718 ();
 FILLCELL_X1 FILLER_0_1_720 ();
 FILLCELL_X1 FILLER_0_1_755 ();
 FILLCELL_X16 FILLER_0_1_776 ();
 FILLCELL_X2 FILLER_0_1_792 ();
 FILLCELL_X1 FILLER_0_1_794 ();
 FILLCELL_X2 FILLER_0_1_815 ();
 FILLCELL_X1 FILLER_0_1_817 ();
 FILLCELL_X1 FILLER_0_1_827 ();
 FILLCELL_X2 FILLER_0_1_837 ();
 FILLCELL_X1 FILLER_0_1_848 ();
 FILLCELL_X1 FILLER_0_1_858 ();
 FILLCELL_X4 FILLER_0_1_869 ();
 FILLCELL_X2 FILLER_0_1_880 ();
 FILLCELL_X2 FILLER_0_1_902 ();
 FILLCELL_X1 FILLER_0_1_934 ();
 FILLCELL_X2 FILLER_0_1_940 ();
 FILLCELL_X2 FILLER_0_1_964 ();
 FILLCELL_X1 FILLER_0_1_986 ();
 FILLCELL_X4 FILLER_0_1_1001 ();
 FILLCELL_X1 FILLER_0_1_1005 ();
 FILLCELL_X1 FILLER_0_1_1031 ();
 FILLCELL_X32 FILLER_0_1_1042 ();
 FILLCELL_X32 FILLER_0_1_1074 ();
 FILLCELL_X32 FILLER_0_1_1106 ();
 FILLCELL_X8 FILLER_0_1_1138 ();
 FILLCELL_X2 FILLER_0_1_1146 ();
 FILLCELL_X32 FILLER_0_2_1 ();
 FILLCELL_X32 FILLER_0_2_33 ();
 FILLCELL_X32 FILLER_0_2_65 ();
 FILLCELL_X32 FILLER_0_2_97 ();
 FILLCELL_X32 FILLER_0_2_129 ();
 FILLCELL_X32 FILLER_0_2_161 ();
 FILLCELL_X32 FILLER_0_2_193 ();
 FILLCELL_X16 FILLER_0_2_225 ();
 FILLCELL_X8 FILLER_0_2_241 ();
 FILLCELL_X4 FILLER_0_2_249 ();
 FILLCELL_X1 FILLER_0_2_258 ();
 FILLCELL_X1 FILLER_0_2_264 ();
 FILLCELL_X1 FILLER_0_2_290 ();
 FILLCELL_X2 FILLER_0_2_301 ();
 FILLCELL_X2 FILLER_0_2_345 ();
 FILLCELL_X1 FILLER_0_2_347 ();
 FILLCELL_X4 FILLER_0_2_383 ();
 FILLCELL_X1 FILLER_0_2_416 ();
 FILLCELL_X2 FILLER_0_2_447 ();
 FILLCELL_X1 FILLER_0_2_449 ();
 FILLCELL_X2 FILLER_0_2_473 ();
 FILLCELL_X2 FILLER_0_2_485 ();
 FILLCELL_X2 FILLER_0_2_497 ();
 FILLCELL_X1 FILLER_0_2_572 ();
 FILLCELL_X4 FILLER_0_2_583 ();
 FILLCELL_X4 FILLER_0_2_617 ();
 FILLCELL_X1 FILLER_0_2_632 ();
 FILLCELL_X4 FILLER_0_2_648 ();
 FILLCELL_X4 FILLER_0_2_659 ();
 FILLCELL_X2 FILLER_0_2_673 ();
 FILLCELL_X1 FILLER_0_2_675 ();
 FILLCELL_X2 FILLER_0_2_757 ();
 FILLCELL_X1 FILLER_0_2_759 ();
 FILLCELL_X1 FILLER_0_2_795 ();
 FILLCELL_X4 FILLER_0_2_815 ();
 FILLCELL_X2 FILLER_0_2_819 ();
 FILLCELL_X4 FILLER_0_2_831 ();
 FILLCELL_X2 FILLER_0_2_835 ();
 FILLCELL_X1 FILLER_0_2_890 ();
 FILLCELL_X1 FILLER_0_2_896 ();
 FILLCELL_X2 FILLER_0_2_966 ();
 FILLCELL_X1 FILLER_0_2_968 ();
 FILLCELL_X1 FILLER_0_2_979 ();
 FILLCELL_X1 FILLER_0_2_990 ();
 FILLCELL_X1 FILLER_0_2_996 ();
 FILLCELL_X1 FILLER_0_2_1007 ();
 FILLCELL_X32 FILLER_0_2_1038 ();
 FILLCELL_X32 FILLER_0_2_1070 ();
 FILLCELL_X32 FILLER_0_2_1102 ();
 FILLCELL_X8 FILLER_0_2_1134 ();
 FILLCELL_X4 FILLER_0_2_1142 ();
 FILLCELL_X2 FILLER_0_2_1146 ();
 FILLCELL_X32 FILLER_0_3_1 ();
 FILLCELL_X32 FILLER_0_3_33 ();
 FILLCELL_X32 FILLER_0_3_65 ();
 FILLCELL_X32 FILLER_0_3_97 ();
 FILLCELL_X32 FILLER_0_3_129 ();
 FILLCELL_X32 FILLER_0_3_161 ();
 FILLCELL_X32 FILLER_0_3_193 ();
 FILLCELL_X8 FILLER_0_3_225 ();
 FILLCELL_X4 FILLER_0_3_233 ();
 FILLCELL_X2 FILLER_0_3_237 ();
 FILLCELL_X4 FILLER_0_3_259 ();
 FILLCELL_X2 FILLER_0_3_330 ();
 FILLCELL_X1 FILLER_0_3_332 ();
 FILLCELL_X1 FILLER_0_3_352 ();
 FILLCELL_X2 FILLER_0_3_363 ();
 FILLCELL_X1 FILLER_0_3_370 ();
 FILLCELL_X1 FILLER_0_3_376 ();
 FILLCELL_X1 FILLER_0_3_392 ();
 FILLCELL_X2 FILLER_0_3_422 ();
 FILLCELL_X1 FILLER_0_3_460 ();
 FILLCELL_X1 FILLER_0_3_485 ();
 FILLCELL_X4 FILLER_0_3_501 ();
 FILLCELL_X4 FILLER_0_3_517 ();
 FILLCELL_X2 FILLER_0_3_531 ();
 FILLCELL_X1 FILLER_0_3_533 ();
 FILLCELL_X1 FILLER_0_3_544 ();
 FILLCELL_X1 FILLER_0_3_555 ();
 FILLCELL_X1 FILLER_0_3_561 ();
 FILLCELL_X1 FILLER_0_3_567 ();
 FILLCELL_X1 FILLER_0_3_578 ();
 FILLCELL_X2 FILLER_0_3_584 ();
 FILLCELL_X2 FILLER_0_3_606 ();
 FILLCELL_X1 FILLER_0_3_608 ();
 FILLCELL_X4 FILLER_0_3_619 ();
 FILLCELL_X2 FILLER_0_3_623 ();
 FILLCELL_X1 FILLER_0_3_625 ();
 FILLCELL_X2 FILLER_0_3_688 ();
 FILLCELL_X1 FILLER_0_3_718 ();
 FILLCELL_X2 FILLER_0_3_733 ();
 FILLCELL_X1 FILLER_0_3_735 ();
 FILLCELL_X8 FILLER_0_3_775 ();
 FILLCELL_X2 FILLER_0_3_853 ();
 FILLCELL_X1 FILLER_0_3_865 ();
 FILLCELL_X1 FILLER_0_3_946 ();
 FILLCELL_X2 FILLER_0_3_954 ();
 FILLCELL_X1 FILLER_0_3_966 ();
 FILLCELL_X1 FILLER_0_3_977 ();
 FILLCELL_X4 FILLER_0_3_992 ();
 FILLCELL_X2 FILLER_0_3_1005 ();
 FILLCELL_X1 FILLER_0_3_1007 ();
 FILLCELL_X2 FILLER_0_3_1027 ();
 FILLCELL_X32 FILLER_0_3_1049 ();
 FILLCELL_X32 FILLER_0_3_1081 ();
 FILLCELL_X32 FILLER_0_3_1113 ();
 FILLCELL_X2 FILLER_0_3_1145 ();
 FILLCELL_X1 FILLER_0_3_1147 ();
 FILLCELL_X32 FILLER_0_4_1 ();
 FILLCELL_X32 FILLER_0_4_33 ();
 FILLCELL_X32 FILLER_0_4_65 ();
 FILLCELL_X32 FILLER_0_4_97 ();
 FILLCELL_X32 FILLER_0_4_129 ();
 FILLCELL_X32 FILLER_0_4_161 ();
 FILLCELL_X32 FILLER_0_4_193 ();
 FILLCELL_X16 FILLER_0_4_225 ();
 FILLCELL_X2 FILLER_0_4_241 ();
 FILLCELL_X2 FILLER_0_4_312 ();
 FILLCELL_X2 FILLER_0_4_355 ();
 FILLCELL_X1 FILLER_0_4_357 ();
 FILLCELL_X4 FILLER_0_4_427 ();
 FILLCELL_X2 FILLER_0_4_441 ();
 FILLCELL_X1 FILLER_0_4_443 ();
 FILLCELL_X1 FILLER_0_4_458 ();
 FILLCELL_X1 FILLER_0_4_469 ();
 FILLCELL_X1 FILLER_0_4_480 ();
 FILLCELL_X4 FILLER_0_4_491 ();
 FILLCELL_X2 FILLER_0_4_519 ();
 FILLCELL_X1 FILLER_0_4_564 ();
 FILLCELL_X8 FILLER_0_4_575 ();
 FILLCELL_X2 FILLER_0_4_583 ();
 FILLCELL_X1 FILLER_0_4_585 ();
 FILLCELL_X16 FILLER_0_4_611 ();
 FILLCELL_X4 FILLER_0_4_627 ();
 FILLCELL_X4 FILLER_0_4_632 ();
 FILLCELL_X1 FILLER_0_4_636 ();
 FILLCELL_X2 FILLER_0_4_647 ();
 FILLCELL_X1 FILLER_0_4_658 ();
 FILLCELL_X16 FILLER_0_4_674 ();
 FILLCELL_X1 FILLER_0_4_700 ();
 FILLCELL_X1 FILLER_0_4_726 ();
 FILLCELL_X2 FILLER_0_4_745 ();
 FILLCELL_X1 FILLER_0_4_747 ();
 FILLCELL_X4 FILLER_0_4_763 ();
 FILLCELL_X1 FILLER_0_4_767 ();
 FILLCELL_X1 FILLER_0_4_788 ();
 FILLCELL_X16 FILLER_0_4_809 ();
 FILLCELL_X1 FILLER_0_4_825 ();
 FILLCELL_X1 FILLER_0_4_842 ();
 FILLCELL_X2 FILLER_0_4_863 ();
 FILLCELL_X1 FILLER_0_4_865 ();
 FILLCELL_X2 FILLER_0_4_940 ();
 FILLCELL_X1 FILLER_0_4_979 ();
 FILLCELL_X4 FILLER_0_4_1005 ();
 FILLCELL_X2 FILLER_0_4_1024 ();
 FILLCELL_X1 FILLER_0_4_1031 ();
 FILLCELL_X1 FILLER_0_4_1036 ();
 FILLCELL_X4 FILLER_0_4_1051 ();
 FILLCELL_X1 FILLER_0_4_1055 ();
 FILLCELL_X32 FILLER_0_4_1066 ();
 FILLCELL_X32 FILLER_0_4_1098 ();
 FILLCELL_X16 FILLER_0_4_1130 ();
 FILLCELL_X2 FILLER_0_4_1146 ();
 FILLCELL_X32 FILLER_0_5_1 ();
 FILLCELL_X32 FILLER_0_5_33 ();
 FILLCELL_X32 FILLER_0_5_65 ();
 FILLCELL_X32 FILLER_0_5_97 ();
 FILLCELL_X32 FILLER_0_5_129 ();
 FILLCELL_X32 FILLER_0_5_161 ();
 FILLCELL_X32 FILLER_0_5_193 ();
 FILLCELL_X4 FILLER_0_5_225 ();
 FILLCELL_X2 FILLER_0_5_254 ();
 FILLCELL_X1 FILLER_0_5_256 ();
 FILLCELL_X1 FILLER_0_5_271 ();
 FILLCELL_X1 FILLER_0_5_282 ();
 FILLCELL_X1 FILLER_0_5_300 ();
 FILLCELL_X4 FILLER_0_5_337 ();
 FILLCELL_X4 FILLER_0_5_351 ();
 FILLCELL_X4 FILLER_0_5_365 ();
 FILLCELL_X1 FILLER_0_5_369 ();
 FILLCELL_X8 FILLER_0_5_389 ();
 FILLCELL_X4 FILLER_0_5_397 ();
 FILLCELL_X1 FILLER_0_5_401 ();
 FILLCELL_X4 FILLER_0_5_432 ();
 FILLCELL_X1 FILLER_0_5_466 ();
 FILLCELL_X4 FILLER_0_5_487 ();
 FILLCELL_X1 FILLER_0_5_518 ();
 FILLCELL_X1 FILLER_0_5_533 ();
 FILLCELL_X2 FILLER_0_5_544 ();
 FILLCELL_X1 FILLER_0_5_546 ();
 FILLCELL_X8 FILLER_0_5_562 ();
 FILLCELL_X2 FILLER_0_5_570 ();
 FILLCELL_X4 FILLER_0_5_604 ();
 FILLCELL_X16 FILLER_0_5_613 ();
 FILLCELL_X2 FILLER_0_5_629 ();
 FILLCELL_X2 FILLER_0_5_646 ();
 FILLCELL_X1 FILLER_0_5_648 ();
 FILLCELL_X4 FILLER_0_5_668 ();
 FILLCELL_X2 FILLER_0_5_687 ();
 FILLCELL_X4 FILLER_0_5_703 ();
 FILLCELL_X1 FILLER_0_5_754 ();
 FILLCELL_X2 FILLER_0_5_770 ();
 FILLCELL_X1 FILLER_0_5_772 ();
 FILLCELL_X1 FILLER_0_5_784 ();
 FILLCELL_X2 FILLER_0_5_800 ();
 FILLCELL_X16 FILLER_0_5_812 ();
 FILLCELL_X1 FILLER_0_5_828 ();
 FILLCELL_X1 FILLER_0_5_858 ();
 FILLCELL_X4 FILLER_0_5_869 ();
 FILLCELL_X2 FILLER_0_5_894 ();
 FILLCELL_X4 FILLER_0_5_906 ();
 FILLCELL_X2 FILLER_0_5_931 ();
 FILLCELL_X1 FILLER_0_5_950 ();
 FILLCELL_X2 FILLER_0_5_998 ();
 FILLCELL_X1 FILLER_0_5_1030 ();
 FILLCELL_X1 FILLER_0_5_1041 ();
 FILLCELL_X32 FILLER_0_5_1057 ();
 FILLCELL_X32 FILLER_0_5_1089 ();
 FILLCELL_X16 FILLER_0_5_1121 ();
 FILLCELL_X8 FILLER_0_5_1137 ();
 FILLCELL_X2 FILLER_0_5_1145 ();
 FILLCELL_X1 FILLER_0_5_1147 ();
 FILLCELL_X32 FILLER_0_6_1 ();
 FILLCELL_X32 FILLER_0_6_33 ();
 FILLCELL_X32 FILLER_0_6_65 ();
 FILLCELL_X32 FILLER_0_6_97 ();
 FILLCELL_X32 FILLER_0_6_129 ();
 FILLCELL_X32 FILLER_0_6_161 ();
 FILLCELL_X16 FILLER_0_6_193 ();
 FILLCELL_X2 FILLER_0_6_209 ();
 FILLCELL_X1 FILLER_0_6_211 ();
 FILLCELL_X2 FILLER_0_6_227 ();
 FILLCELL_X1 FILLER_0_6_229 ();
 FILLCELL_X2 FILLER_0_6_277 ();
 FILLCELL_X1 FILLER_0_6_289 ();
 FILLCELL_X1 FILLER_0_6_305 ();
 FILLCELL_X2 FILLER_0_6_325 ();
 FILLCELL_X1 FILLER_0_6_327 ();
 FILLCELL_X8 FILLER_0_6_362 ();
 FILLCELL_X16 FILLER_0_6_379 ();
 FILLCELL_X8 FILLER_0_6_395 ();
 FILLCELL_X4 FILLER_0_6_403 ();
 FILLCELL_X1 FILLER_0_6_407 ();
 FILLCELL_X1 FILLER_0_6_437 ();
 FILLCELL_X1 FILLER_0_6_448 ();
 FILLCELL_X4 FILLER_0_6_464 ();
 FILLCELL_X2 FILLER_0_6_475 ();
 FILLCELL_X1 FILLER_0_6_497 ();
 FILLCELL_X2 FILLER_0_6_518 ();
 FILLCELL_X2 FILLER_0_6_540 ();
 FILLCELL_X2 FILLER_0_6_556 ();
 FILLCELL_X8 FILLER_0_6_568 ();
 FILLCELL_X2 FILLER_0_6_576 ();
 FILLCELL_X1 FILLER_0_6_603 ();
 FILLCELL_X16 FILLER_0_6_614 ();
 FILLCELL_X1 FILLER_0_6_630 ();
 FILLCELL_X8 FILLER_0_6_632 ();
 FILLCELL_X2 FILLER_0_6_640 ();
 FILLCELL_X1 FILLER_0_6_642 ();
 FILLCELL_X1 FILLER_0_6_658 ();
 FILLCELL_X4 FILLER_0_6_699 ();
 FILLCELL_X1 FILLER_0_6_750 ();
 FILLCELL_X2 FILLER_0_6_776 ();
 FILLCELL_X4 FILLER_0_6_788 ();
 FILLCELL_X16 FILLER_0_6_802 ();
 FILLCELL_X4 FILLER_0_6_818 ();
 FILLCELL_X2 FILLER_0_6_822 ();
 FILLCELL_X1 FILLER_0_6_824 ();
 FILLCELL_X1 FILLER_0_6_872 ();
 FILLCELL_X1 FILLER_0_6_880 ();
 FILLCELL_X1 FILLER_0_6_924 ();
 FILLCELL_X1 FILLER_0_6_940 ();
 FILLCELL_X2 FILLER_0_6_982 ();
 FILLCELL_X4 FILLER_0_6_1010 ();
 FILLCELL_X1 FILLER_0_6_1044 ();
 FILLCELL_X32 FILLER_0_6_1055 ();
 FILLCELL_X32 FILLER_0_6_1087 ();
 FILLCELL_X16 FILLER_0_6_1119 ();
 FILLCELL_X8 FILLER_0_6_1135 ();
 FILLCELL_X4 FILLER_0_6_1143 ();
 FILLCELL_X1 FILLER_0_6_1147 ();
 FILLCELL_X32 FILLER_0_7_1 ();
 FILLCELL_X32 FILLER_0_7_33 ();
 FILLCELL_X32 FILLER_0_7_65 ();
 FILLCELL_X32 FILLER_0_7_97 ();
 FILLCELL_X32 FILLER_0_7_129 ();
 FILLCELL_X32 FILLER_0_7_161 ();
 FILLCELL_X8 FILLER_0_7_193 ();
 FILLCELL_X2 FILLER_0_7_201 ();
 FILLCELL_X1 FILLER_0_7_203 ();
 FILLCELL_X1 FILLER_0_7_219 ();
 FILLCELL_X2 FILLER_0_7_238 ();
 FILLCELL_X1 FILLER_0_7_240 ();
 FILLCELL_X1 FILLER_0_7_306 ();
 FILLCELL_X2 FILLER_0_7_317 ();
 FILLCELL_X1 FILLER_0_7_319 ();
 FILLCELL_X8 FILLER_0_7_377 ();
 FILLCELL_X2 FILLER_0_7_385 ();
 FILLCELL_X2 FILLER_0_7_397 ();
 FILLCELL_X1 FILLER_0_7_436 ();
 FILLCELL_X1 FILLER_0_7_510 ();
 FILLCELL_X1 FILLER_0_7_526 ();
 FILLCELL_X2 FILLER_0_7_569 ();
 FILLCELL_X1 FILLER_0_7_581 ();
 FILLCELL_X4 FILLER_0_7_596 ();
 FILLCELL_X2 FILLER_0_7_600 ();
 FILLCELL_X1 FILLER_0_7_602 ();
 FILLCELL_X16 FILLER_0_7_613 ();
 FILLCELL_X8 FILLER_0_7_629 ();
 FILLCELL_X4 FILLER_0_7_637 ();
 FILLCELL_X4 FILLER_0_7_661 ();
 FILLCELL_X2 FILLER_0_7_675 ();
 FILLCELL_X1 FILLER_0_7_677 ();
 FILLCELL_X1 FILLER_0_7_709 ();
 FILLCELL_X2 FILLER_0_7_752 ();
 FILLCELL_X1 FILLER_0_7_754 ();
 FILLCELL_X8 FILLER_0_7_809 ();
 FILLCELL_X4 FILLER_0_7_817 ();
 FILLCELL_X1 FILLER_0_7_831 ();
 FILLCELL_X1 FILLER_0_7_866 ();
 FILLCELL_X4 FILLER_0_7_884 ();
 FILLCELL_X2 FILLER_0_7_915 ();
 FILLCELL_X1 FILLER_0_7_917 ();
 FILLCELL_X1 FILLER_0_7_935 ();
 FILLCELL_X2 FILLER_0_7_993 ();
 FILLCELL_X2 FILLER_0_7_1005 ();
 FILLCELL_X1 FILLER_0_7_1007 ();
 FILLCELL_X2 FILLER_0_7_1018 ();
 FILLCELL_X1 FILLER_0_7_1020 ();
 FILLCELL_X2 FILLER_0_7_1026 ();
 FILLCELL_X1 FILLER_0_7_1028 ();
 FILLCELL_X32 FILLER_0_7_1039 ();
 FILLCELL_X32 FILLER_0_7_1071 ();
 FILLCELL_X32 FILLER_0_7_1103 ();
 FILLCELL_X8 FILLER_0_7_1135 ();
 FILLCELL_X4 FILLER_0_7_1143 ();
 FILLCELL_X1 FILLER_0_7_1147 ();
 FILLCELL_X32 FILLER_0_8_1 ();
 FILLCELL_X32 FILLER_0_8_33 ();
 FILLCELL_X32 FILLER_0_8_65 ();
 FILLCELL_X32 FILLER_0_8_97 ();
 FILLCELL_X32 FILLER_0_8_129 ();
 FILLCELL_X32 FILLER_0_8_161 ();
 FILLCELL_X16 FILLER_0_8_193 ();
 FILLCELL_X4 FILLER_0_8_209 ();
 FILLCELL_X1 FILLER_0_8_263 ();
 FILLCELL_X4 FILLER_0_8_288 ();
 FILLCELL_X8 FILLER_0_8_374 ();
 FILLCELL_X1 FILLER_0_8_382 ();
 FILLCELL_X2 FILLER_0_8_429 ();
 FILLCELL_X1 FILLER_0_8_438 ();
 FILLCELL_X1 FILLER_0_8_511 ();
 FILLCELL_X1 FILLER_0_8_522 ();
 FILLCELL_X2 FILLER_0_8_569 ();
 FILLCELL_X2 FILLER_0_8_586 ();
 FILLCELL_X1 FILLER_0_8_588 ();
 FILLCELL_X8 FILLER_0_8_603 ();
 FILLCELL_X4 FILLER_0_8_611 ();
 FILLCELL_X1 FILLER_0_8_615 ();
 FILLCELL_X2 FILLER_0_8_664 ();
 FILLCELL_X1 FILLER_0_8_666 ();
 FILLCELL_X2 FILLER_0_8_684 ();
 FILLCELL_X1 FILLER_0_8_686 ();
 FILLCELL_X2 FILLER_0_8_743 ();
 FILLCELL_X1 FILLER_0_8_770 ();
 FILLCELL_X2 FILLER_0_8_787 ();
 FILLCELL_X1 FILLER_0_8_789 ();
 FILLCELL_X4 FILLER_0_8_805 ();
 FILLCELL_X2 FILLER_0_8_809 ();
 FILLCELL_X1 FILLER_0_8_811 ();
 FILLCELL_X1 FILLER_0_8_900 ();
 FILLCELL_X2 FILLER_0_8_908 ();
 FILLCELL_X1 FILLER_0_8_941 ();
 FILLCELL_X2 FILLER_0_8_959 ();
 FILLCELL_X4 FILLER_0_8_984 ();
 FILLCELL_X1 FILLER_0_8_998 ();
 FILLCELL_X1 FILLER_0_8_1009 ();
 FILLCELL_X1 FILLER_0_8_1020 ();
 FILLCELL_X1 FILLER_0_8_1030 ();
 FILLCELL_X1 FILLER_0_8_1041 ();
 FILLCELL_X32 FILLER_0_8_1052 ();
 FILLCELL_X32 FILLER_0_8_1084 ();
 FILLCELL_X32 FILLER_0_8_1116 ();
 FILLCELL_X32 FILLER_0_9_1 ();
 FILLCELL_X32 FILLER_0_9_33 ();
 FILLCELL_X32 FILLER_0_9_65 ();
 FILLCELL_X32 FILLER_0_9_97 ();
 FILLCELL_X32 FILLER_0_9_129 ();
 FILLCELL_X32 FILLER_0_9_161 ();
 FILLCELL_X16 FILLER_0_9_193 ();
 FILLCELL_X2 FILLER_0_9_209 ();
 FILLCELL_X2 FILLER_0_9_221 ();
 FILLCELL_X1 FILLER_0_9_242 ();
 FILLCELL_X2 FILLER_0_9_253 ();
 FILLCELL_X2 FILLER_0_9_280 ();
 FILLCELL_X1 FILLER_0_9_282 ();
 FILLCELL_X2 FILLER_0_9_371 ();
 FILLCELL_X1 FILLER_0_9_388 ();
 FILLCELL_X1 FILLER_0_9_394 ();
 FILLCELL_X1 FILLER_0_9_400 ();
 FILLCELL_X4 FILLER_0_9_411 ();
 FILLCELL_X2 FILLER_0_9_425 ();
 FILLCELL_X2 FILLER_0_9_475 ();
 FILLCELL_X1 FILLER_0_9_477 ();
 FILLCELL_X1 FILLER_0_9_495 ();
 FILLCELL_X4 FILLER_0_9_530 ();
 FILLCELL_X1 FILLER_0_9_544 ();
 FILLCELL_X2 FILLER_0_9_572 ();
 FILLCELL_X1 FILLER_0_9_574 ();
 FILLCELL_X8 FILLER_0_9_585 ();
 FILLCELL_X4 FILLER_0_9_593 ();
 FILLCELL_X1 FILLER_0_9_597 ();
 FILLCELL_X2 FILLER_0_9_603 ();
 FILLCELL_X4 FILLER_0_9_615 ();
 FILLCELL_X2 FILLER_0_9_619 ();
 FILLCELL_X2 FILLER_0_9_626 ();
 FILLCELL_X1 FILLER_0_9_702 ();
 FILLCELL_X1 FILLER_0_9_747 ();
 FILLCELL_X1 FILLER_0_9_763 ();
 FILLCELL_X1 FILLER_0_9_773 ();
 FILLCELL_X2 FILLER_0_9_800 ();
 FILLCELL_X4 FILLER_0_9_812 ();
 FILLCELL_X2 FILLER_0_9_816 ();
 FILLCELL_X1 FILLER_0_9_818 ();
 FILLCELL_X2 FILLER_0_9_834 ();
 FILLCELL_X1 FILLER_0_9_843 ();
 FILLCELL_X2 FILLER_0_9_869 ();
 FILLCELL_X1 FILLER_0_9_900 ();
 FILLCELL_X1 FILLER_0_9_936 ();
 FILLCELL_X1 FILLER_0_9_946 ();
 FILLCELL_X1 FILLER_0_9_954 ();
 FILLCELL_X4 FILLER_0_9_1007 ();
 FILLCELL_X2 FILLER_0_9_1035 ();
 FILLCELL_X32 FILLER_0_9_1057 ();
 FILLCELL_X32 FILLER_0_9_1089 ();
 FILLCELL_X16 FILLER_0_9_1121 ();
 FILLCELL_X8 FILLER_0_9_1137 ();
 FILLCELL_X2 FILLER_0_9_1145 ();
 FILLCELL_X1 FILLER_0_9_1147 ();
 FILLCELL_X32 FILLER_0_10_1 ();
 FILLCELL_X32 FILLER_0_10_33 ();
 FILLCELL_X32 FILLER_0_10_65 ();
 FILLCELL_X32 FILLER_0_10_97 ();
 FILLCELL_X32 FILLER_0_10_129 ();
 FILLCELL_X32 FILLER_0_10_161 ();
 FILLCELL_X8 FILLER_0_10_193 ();
 FILLCELL_X1 FILLER_0_10_221 ();
 FILLCELL_X1 FILLER_0_10_271 ();
 FILLCELL_X2 FILLER_0_10_299 ();
 FILLCELL_X1 FILLER_0_10_301 ();
 FILLCELL_X1 FILLER_0_10_327 ();
 FILLCELL_X1 FILLER_0_10_337 ();
 FILLCELL_X1 FILLER_0_10_357 ();
 FILLCELL_X4 FILLER_0_10_377 ();
 FILLCELL_X1 FILLER_0_10_391 ();
 FILLCELL_X8 FILLER_0_10_396 ();
 FILLCELL_X4 FILLER_0_10_404 ();
 FILLCELL_X2 FILLER_0_10_408 ();
 FILLCELL_X1 FILLER_0_10_410 ();
 FILLCELL_X2 FILLER_0_10_443 ();
 FILLCELL_X4 FILLER_0_10_455 ();
 FILLCELL_X2 FILLER_0_10_525 ();
 FILLCELL_X8 FILLER_0_10_581 ();
 FILLCELL_X4 FILLER_0_10_589 ();
 FILLCELL_X2 FILLER_0_10_593 ();
 FILLCELL_X1 FILLER_0_10_595 ();
 FILLCELL_X8 FILLER_0_10_606 ();
 FILLCELL_X4 FILLER_0_10_614 ();
 FILLCELL_X2 FILLER_0_10_618 ();
 FILLCELL_X1 FILLER_0_10_620 ();
 FILLCELL_X2 FILLER_0_10_632 ();
 FILLCELL_X1 FILLER_0_10_644 ();
 FILLCELL_X2 FILLER_0_10_662 ();
 FILLCELL_X1 FILLER_0_10_714 ();
 FILLCELL_X2 FILLER_0_10_755 ();
 FILLCELL_X1 FILLER_0_10_789 ();
 FILLCELL_X16 FILLER_0_10_805 ();
 FILLCELL_X1 FILLER_0_10_834 ();
 FILLCELL_X4 FILLER_0_10_852 ();
 FILLCELL_X2 FILLER_0_10_866 ();
 FILLCELL_X1 FILLER_0_10_868 ();
 FILLCELL_X2 FILLER_0_10_906 ();
 FILLCELL_X1 FILLER_0_10_908 ();
 FILLCELL_X1 FILLER_0_10_946 ();
 FILLCELL_X4 FILLER_0_10_982 ();
 FILLCELL_X2 FILLER_0_10_1006 ();
 FILLCELL_X1 FILLER_0_10_1008 ();
 FILLCELL_X1 FILLER_0_10_1052 ();
 FILLCELL_X32 FILLER_0_10_1063 ();
 FILLCELL_X32 FILLER_0_10_1095 ();
 FILLCELL_X16 FILLER_0_10_1127 ();
 FILLCELL_X4 FILLER_0_10_1143 ();
 FILLCELL_X1 FILLER_0_10_1147 ();
 FILLCELL_X32 FILLER_0_11_1 ();
 FILLCELL_X32 FILLER_0_11_33 ();
 FILLCELL_X32 FILLER_0_11_65 ();
 FILLCELL_X32 FILLER_0_11_97 ();
 FILLCELL_X32 FILLER_0_11_129 ();
 FILLCELL_X32 FILLER_0_11_161 ();
 FILLCELL_X8 FILLER_0_11_193 ();
 FILLCELL_X2 FILLER_0_11_211 ();
 FILLCELL_X1 FILLER_0_11_213 ();
 FILLCELL_X1 FILLER_0_11_268 ();
 FILLCELL_X1 FILLER_0_11_322 ();
 FILLCELL_X1 FILLER_0_11_361 ();
 FILLCELL_X2 FILLER_0_11_415 ();
 FILLCELL_X1 FILLER_0_11_417 ();
 FILLCELL_X1 FILLER_0_11_487 ();
 FILLCELL_X1 FILLER_0_11_520 ();
 FILLCELL_X2 FILLER_0_11_583 ();
 FILLCELL_X1 FILLER_0_11_585 ();
 FILLCELL_X16 FILLER_0_11_606 ();
 FILLCELL_X8 FILLER_0_11_622 ();
 FILLCELL_X4 FILLER_0_11_630 ();
 FILLCELL_X1 FILLER_0_11_634 ();
 FILLCELL_X4 FILLER_0_11_655 ();
 FILLCELL_X1 FILLER_0_11_659 ();
 FILLCELL_X2 FILLER_0_11_760 ();
 FILLCELL_X1 FILLER_0_11_762 ();
 FILLCELL_X1 FILLER_0_11_785 ();
 FILLCELL_X16 FILLER_0_11_802 ();
 FILLCELL_X8 FILLER_0_11_818 ();
 FILLCELL_X4 FILLER_0_11_836 ();
 FILLCELL_X2 FILLER_0_11_840 ();
 FILLCELL_X1 FILLER_0_11_842 ();
 FILLCELL_X1 FILLER_0_11_860 ();
 FILLCELL_X1 FILLER_0_11_880 ();
 FILLCELL_X4 FILLER_0_11_903 ();
 FILLCELL_X1 FILLER_0_11_992 ();
 FILLCELL_X1 FILLER_0_11_1041 ();
 FILLCELL_X32 FILLER_0_11_1057 ();
 FILLCELL_X32 FILLER_0_11_1089 ();
 FILLCELL_X16 FILLER_0_11_1121 ();
 FILLCELL_X8 FILLER_0_11_1137 ();
 FILLCELL_X2 FILLER_0_11_1145 ();
 FILLCELL_X1 FILLER_0_11_1147 ();
 FILLCELL_X32 FILLER_0_12_1 ();
 FILLCELL_X32 FILLER_0_12_33 ();
 FILLCELL_X32 FILLER_0_12_65 ();
 FILLCELL_X32 FILLER_0_12_97 ();
 FILLCELL_X32 FILLER_0_12_129 ();
 FILLCELL_X32 FILLER_0_12_161 ();
 FILLCELL_X1 FILLER_0_12_193 ();
 FILLCELL_X2 FILLER_0_12_228 ();
 FILLCELL_X1 FILLER_0_12_267 ();
 FILLCELL_X4 FILLER_0_12_278 ();
 FILLCELL_X2 FILLER_0_12_307 ();
 FILLCELL_X1 FILLER_0_12_309 ();
 FILLCELL_X1 FILLER_0_12_319 ();
 FILLCELL_X4 FILLER_0_12_423 ();
 FILLCELL_X2 FILLER_0_12_471 ();
 FILLCELL_X1 FILLER_0_12_473 ();
 FILLCELL_X2 FILLER_0_12_491 ();
 FILLCELL_X1 FILLER_0_12_493 ();
 FILLCELL_X1 FILLER_0_12_510 ();
 FILLCELL_X1 FILLER_0_12_533 ();
 FILLCELL_X2 FILLER_0_12_580 ();
 FILLCELL_X2 FILLER_0_12_587 ();
 FILLCELL_X1 FILLER_0_12_594 ();
 FILLCELL_X16 FILLER_0_12_605 ();
 FILLCELL_X1 FILLER_0_12_632 ();
 FILLCELL_X4 FILLER_0_12_643 ();
 FILLCELL_X1 FILLER_0_12_647 ();
 FILLCELL_X4 FILLER_0_12_683 ();
 FILLCELL_X2 FILLER_0_12_734 ();
 FILLCELL_X4 FILLER_0_12_813 ();
 FILLCELL_X2 FILLER_0_12_817 ();
 FILLCELL_X8 FILLER_0_12_824 ();
 FILLCELL_X4 FILLER_0_12_832 ();
 FILLCELL_X1 FILLER_0_12_836 ();
 FILLCELL_X2 FILLER_0_12_856 ();
 FILLCELL_X1 FILLER_0_12_858 ();
 FILLCELL_X1 FILLER_0_12_869 ();
 FILLCELL_X2 FILLER_0_12_894 ();
 FILLCELL_X1 FILLER_0_12_896 ();
 FILLCELL_X1 FILLER_0_12_936 ();
 FILLCELL_X2 FILLER_0_12_1018 ();
 FILLCELL_X2 FILLER_0_12_1030 ();
 FILLCELL_X1 FILLER_0_12_1041 ();
 FILLCELL_X32 FILLER_0_12_1052 ();
 FILLCELL_X32 FILLER_0_12_1084 ();
 FILLCELL_X32 FILLER_0_12_1116 ();
 FILLCELL_X32 FILLER_0_13_1 ();
 FILLCELL_X32 FILLER_0_13_33 ();
 FILLCELL_X32 FILLER_0_13_65 ();
 FILLCELL_X32 FILLER_0_13_97 ();
 FILLCELL_X32 FILLER_0_13_129 ();
 FILLCELL_X16 FILLER_0_13_161 ();
 FILLCELL_X8 FILLER_0_13_177 ();
 FILLCELL_X4 FILLER_0_13_185 ();
 FILLCELL_X2 FILLER_0_13_189 ();
 FILLCELL_X1 FILLER_0_13_191 ();
 FILLCELL_X2 FILLER_0_13_216 ();
 FILLCELL_X2 FILLER_0_13_228 ();
 FILLCELL_X1 FILLER_0_13_230 ();
 FILLCELL_X2 FILLER_0_13_241 ();
 FILLCELL_X1 FILLER_0_13_243 ();
 FILLCELL_X1 FILLER_0_13_254 ();
 FILLCELL_X2 FILLER_0_13_342 ();
 FILLCELL_X2 FILLER_0_13_354 ();
 FILLCELL_X1 FILLER_0_13_356 ();
 FILLCELL_X1 FILLER_0_13_408 ();
 FILLCELL_X4 FILLER_0_13_415 ();
 FILLCELL_X2 FILLER_0_13_419 ();
 FILLCELL_X1 FILLER_0_13_421 ();
 FILLCELL_X1 FILLER_0_13_439 ();
 FILLCELL_X1 FILLER_0_13_464 ();
 FILLCELL_X2 FILLER_0_13_504 ();
 FILLCELL_X1 FILLER_0_13_551 ();
 FILLCELL_X4 FILLER_0_13_593 ();
 FILLCELL_X8 FILLER_0_13_612 ();
 FILLCELL_X4 FILLER_0_13_620 ();
 FILLCELL_X2 FILLER_0_13_624 ();
 FILLCELL_X1 FILLER_0_13_635 ();
 FILLCELL_X1 FILLER_0_13_651 ();
 FILLCELL_X2 FILLER_0_13_659 ();
 FILLCELL_X4 FILLER_0_13_710 ();
 FILLCELL_X2 FILLER_0_13_752 ();
 FILLCELL_X2 FILLER_0_13_764 ();
 FILLCELL_X1 FILLER_0_13_803 ();
 FILLCELL_X2 FILLER_0_13_821 ();
 FILLCELL_X1 FILLER_0_13_823 ();
 FILLCELL_X4 FILLER_0_13_849 ();
 FILLCELL_X1 FILLER_0_13_860 ();
 FILLCELL_X1 FILLER_0_13_924 ();
 FILLCELL_X1 FILLER_0_13_975 ();
 FILLCELL_X1 FILLER_0_13_1003 ();
 FILLCELL_X2 FILLER_0_13_1013 ();
 FILLCELL_X32 FILLER_0_13_1039 ();
 FILLCELL_X32 FILLER_0_13_1071 ();
 FILLCELL_X32 FILLER_0_13_1103 ();
 FILLCELL_X8 FILLER_0_13_1135 ();
 FILLCELL_X4 FILLER_0_13_1143 ();
 FILLCELL_X1 FILLER_0_13_1147 ();
 FILLCELL_X32 FILLER_0_14_1 ();
 FILLCELL_X32 FILLER_0_14_33 ();
 FILLCELL_X32 FILLER_0_14_65 ();
 FILLCELL_X32 FILLER_0_14_97 ();
 FILLCELL_X32 FILLER_0_14_129 ();
 FILLCELL_X32 FILLER_0_14_161 ();
 FILLCELL_X4 FILLER_0_14_193 ();
 FILLCELL_X4 FILLER_0_14_214 ();
 FILLCELL_X1 FILLER_0_14_227 ();
 FILLCELL_X2 FILLER_0_14_252 ();
 FILLCELL_X1 FILLER_0_14_301 ();
 FILLCELL_X2 FILLER_0_14_317 ();
 FILLCELL_X1 FILLER_0_14_319 ();
 FILLCELL_X2 FILLER_0_14_358 ();
 FILLCELL_X2 FILLER_0_14_384 ();
 FILLCELL_X2 FILLER_0_14_396 ();
 FILLCELL_X2 FILLER_0_14_408 ();
 FILLCELL_X4 FILLER_0_14_416 ();
 FILLCELL_X2 FILLER_0_14_420 ();
 FILLCELL_X2 FILLER_0_14_432 ();
 FILLCELL_X2 FILLER_0_14_451 ();
 FILLCELL_X1 FILLER_0_14_453 ();
 FILLCELL_X2 FILLER_0_14_471 ();
 FILLCELL_X1 FILLER_0_14_507 ();
 FILLCELL_X1 FILLER_0_14_515 ();
 FILLCELL_X1 FILLER_0_14_562 ();
 FILLCELL_X2 FILLER_0_14_570 ();
 FILLCELL_X8 FILLER_0_14_587 ();
 FILLCELL_X4 FILLER_0_14_605 ();
 FILLCELL_X2 FILLER_0_14_609 ();
 FILLCELL_X4 FILLER_0_14_626 ();
 FILLCELL_X1 FILLER_0_14_630 ();
 FILLCELL_X1 FILLER_0_14_637 ();
 FILLCELL_X2 FILLER_0_14_676 ();
 FILLCELL_X1 FILLER_0_14_678 ();
 FILLCELL_X2 FILLER_0_14_709 ();
 FILLCELL_X4 FILLER_0_14_720 ();
 FILLCELL_X2 FILLER_0_14_761 ();
 FILLCELL_X4 FILLER_0_14_790 ();
 FILLCELL_X1 FILLER_0_14_804 ();
 FILLCELL_X2 FILLER_0_14_812 ();
 FILLCELL_X1 FILLER_0_14_864 ();
 FILLCELL_X4 FILLER_0_14_898 ();
 FILLCELL_X4 FILLER_0_14_919 ();
 FILLCELL_X1 FILLER_0_14_961 ();
 FILLCELL_X2 FILLER_0_14_983 ();
 FILLCELL_X32 FILLER_0_14_1052 ();
 FILLCELL_X32 FILLER_0_14_1084 ();
 FILLCELL_X32 FILLER_0_14_1116 ();
 FILLCELL_X32 FILLER_0_15_1 ();
 FILLCELL_X32 FILLER_0_15_33 ();
 FILLCELL_X32 FILLER_0_15_65 ();
 FILLCELL_X32 FILLER_0_15_97 ();
 FILLCELL_X32 FILLER_0_15_129 ();
 FILLCELL_X32 FILLER_0_15_161 ();
 FILLCELL_X8 FILLER_0_15_193 ();
 FILLCELL_X1 FILLER_0_15_201 ();
 FILLCELL_X1 FILLER_0_15_229 ();
 FILLCELL_X2 FILLER_0_15_277 ();
 FILLCELL_X1 FILLER_0_15_279 ();
 FILLCELL_X2 FILLER_0_15_315 ();
 FILLCELL_X1 FILLER_0_15_355 ();
 FILLCELL_X2 FILLER_0_15_377 ();
 FILLCELL_X1 FILLER_0_15_379 ();
 FILLCELL_X1 FILLER_0_15_390 ();
 FILLCELL_X4 FILLER_0_15_407 ();
 FILLCELL_X4 FILLER_0_15_430 ();
 FILLCELL_X2 FILLER_0_15_439 ();
 FILLCELL_X1 FILLER_0_15_441 ();
 FILLCELL_X2 FILLER_0_15_481 ();
 FILLCELL_X1 FILLER_0_15_483 ();
 FILLCELL_X2 FILLER_0_15_515 ();
 FILLCELL_X2 FILLER_0_15_527 ();
 FILLCELL_X1 FILLER_0_15_529 ();
 FILLCELL_X2 FILLER_0_15_540 ();
 FILLCELL_X1 FILLER_0_15_549 ();
 FILLCELL_X16 FILLER_0_15_591 ();
 FILLCELL_X4 FILLER_0_15_607 ();
 FILLCELL_X2 FILLER_0_15_647 ();
 FILLCELL_X1 FILLER_0_15_649 ();
 FILLCELL_X2 FILLER_0_15_677 ();
 FILLCELL_X1 FILLER_0_15_679 ();
 FILLCELL_X4 FILLER_0_15_755 ();
 FILLCELL_X2 FILLER_0_15_809 ();
 FILLCELL_X1 FILLER_0_15_818 ();
 FILLCELL_X8 FILLER_0_15_826 ();
 FILLCELL_X1 FILLER_0_15_848 ();
 FILLCELL_X1 FILLER_0_15_863 ();
 FILLCELL_X2 FILLER_0_15_881 ();
 FILLCELL_X8 FILLER_0_15_906 ();
 FILLCELL_X4 FILLER_0_15_921 ();
 FILLCELL_X2 FILLER_0_15_925 ();
 FILLCELL_X2 FILLER_0_15_956 ();
 FILLCELL_X1 FILLER_0_15_975 ();
 FILLCELL_X2 FILLER_0_15_986 ();
 FILLCELL_X2 FILLER_0_15_998 ();
 FILLCELL_X4 FILLER_0_15_1009 ();
 FILLCELL_X4 FILLER_0_15_1018 ();
 FILLCELL_X2 FILLER_0_15_1022 ();
 FILLCELL_X1 FILLER_0_15_1024 ();
 FILLCELL_X4 FILLER_0_15_1044 ();
 FILLCELL_X1 FILLER_0_15_1048 ();
 FILLCELL_X32 FILLER_0_15_1059 ();
 FILLCELL_X32 FILLER_0_15_1091 ();
 FILLCELL_X16 FILLER_0_15_1123 ();
 FILLCELL_X8 FILLER_0_15_1139 ();
 FILLCELL_X1 FILLER_0_15_1147 ();
 FILLCELL_X32 FILLER_0_16_1 ();
 FILLCELL_X32 FILLER_0_16_33 ();
 FILLCELL_X32 FILLER_0_16_65 ();
 FILLCELL_X32 FILLER_0_16_97 ();
 FILLCELL_X32 FILLER_0_16_129 ();
 FILLCELL_X32 FILLER_0_16_161 ();
 FILLCELL_X4 FILLER_0_16_193 ();
 FILLCELL_X2 FILLER_0_16_197 ();
 FILLCELL_X1 FILLER_0_16_227 ();
 FILLCELL_X2 FILLER_0_16_255 ();
 FILLCELL_X2 FILLER_0_16_284 ();
 FILLCELL_X2 FILLER_0_16_295 ();
 FILLCELL_X1 FILLER_0_16_297 ();
 FILLCELL_X2 FILLER_0_16_363 ();
 FILLCELL_X1 FILLER_0_16_384 ();
 FILLCELL_X16 FILLER_0_16_403 ();
 FILLCELL_X8 FILLER_0_16_419 ();
 FILLCELL_X2 FILLER_0_16_427 ();
 FILLCELL_X1 FILLER_0_16_429 ();
 FILLCELL_X2 FILLER_0_16_443 ();
 FILLCELL_X4 FILLER_0_16_460 ();
 FILLCELL_X1 FILLER_0_16_488 ();
 FILLCELL_X2 FILLER_0_16_526 ();
 FILLCELL_X2 FILLER_0_16_571 ();
 FILLCELL_X1 FILLER_0_16_573 ();
 FILLCELL_X2 FILLER_0_16_589 ();
 FILLCELL_X1 FILLER_0_16_591 ();
 FILLCELL_X8 FILLER_0_16_604 ();
 FILLCELL_X2 FILLER_0_16_612 ();
 FILLCELL_X1 FILLER_0_16_614 ();
 FILLCELL_X1 FILLER_0_16_618 ();
 FILLCELL_X1 FILLER_0_16_630 ();
 FILLCELL_X4 FILLER_0_16_642 ();
 FILLCELL_X1 FILLER_0_16_646 ();
 FILLCELL_X1 FILLER_0_16_674 ();
 FILLCELL_X1 FILLER_0_16_731 ();
 FILLCELL_X4 FILLER_0_16_806 ();
 FILLCELL_X1 FILLER_0_16_810 ();
 FILLCELL_X8 FILLER_0_16_835 ();
 FILLCELL_X4 FILLER_0_16_853 ();
 FILLCELL_X2 FILLER_0_16_857 ();
 FILLCELL_X1 FILLER_0_16_859 ();
 FILLCELL_X2 FILLER_0_16_864 ();
 FILLCELL_X1 FILLER_0_16_866 ();
 FILLCELL_X1 FILLER_0_16_890 ();
 FILLCELL_X4 FILLER_0_16_899 ();
 FILLCELL_X2 FILLER_0_16_975 ();
 FILLCELL_X1 FILLER_0_16_977 ();
 FILLCELL_X2 FILLER_0_16_995 ();
 FILLCELL_X1 FILLER_0_16_997 ();
 FILLCELL_X2 FILLER_0_16_1008 ();
 FILLCELL_X1 FILLER_0_16_1010 ();
 FILLCELL_X2 FILLER_0_16_1021 ();
 FILLCELL_X1 FILLER_0_16_1023 ();
 FILLCELL_X2 FILLER_0_16_1043 ();
 FILLCELL_X2 FILLER_0_16_1050 ();
 FILLCELL_X1 FILLER_0_16_1052 ();
 FILLCELL_X32 FILLER_0_16_1068 ();
 FILLCELL_X32 FILLER_0_16_1100 ();
 FILLCELL_X16 FILLER_0_16_1132 ();
 FILLCELL_X32 FILLER_0_17_1 ();
 FILLCELL_X32 FILLER_0_17_33 ();
 FILLCELL_X32 FILLER_0_17_65 ();
 FILLCELL_X32 FILLER_0_17_97 ();
 FILLCELL_X32 FILLER_0_17_129 ();
 FILLCELL_X32 FILLER_0_17_161 ();
 FILLCELL_X16 FILLER_0_17_193 ();
 FILLCELL_X1 FILLER_0_17_209 ();
 FILLCELL_X2 FILLER_0_17_230 ();
 FILLCELL_X2 FILLER_0_17_263 ();
 FILLCELL_X1 FILLER_0_17_275 ();
 FILLCELL_X1 FILLER_0_17_294 ();
 FILLCELL_X1 FILLER_0_17_322 ();
 FILLCELL_X1 FILLER_0_17_333 ();
 FILLCELL_X2 FILLER_0_17_362 ();
 FILLCELL_X2 FILLER_0_17_417 ();
 FILLCELL_X2 FILLER_0_17_460 ();
 FILLCELL_X2 FILLER_0_17_472 ();
 FILLCELL_X1 FILLER_0_17_488 ();
 FILLCELL_X2 FILLER_0_17_540 ();
 FILLCELL_X1 FILLER_0_17_559 ();
 FILLCELL_X1 FILLER_0_17_570 ();
 FILLCELL_X1 FILLER_0_17_581 ();
 FILLCELL_X2 FILLER_0_17_592 ();
 FILLCELL_X1 FILLER_0_17_594 ();
 FILLCELL_X1 FILLER_0_17_600 ();
 FILLCELL_X2 FILLER_0_17_632 ();
 FILLCELL_X1 FILLER_0_17_719 ();
 FILLCELL_X2 FILLER_0_17_730 ();
 FILLCELL_X1 FILLER_0_17_742 ();
 FILLCELL_X2 FILLER_0_17_763 ();
 FILLCELL_X1 FILLER_0_17_765 ();
 FILLCELL_X1 FILLER_0_17_787 ();
 FILLCELL_X2 FILLER_0_17_826 ();
 FILLCELL_X1 FILLER_0_17_863 ();
 FILLCELL_X1 FILLER_0_17_877 ();
 FILLCELL_X1 FILLER_0_17_882 ();
 FILLCELL_X2 FILLER_0_17_893 ();
 FILLCELL_X2 FILLER_0_17_920 ();
 FILLCELL_X4 FILLER_0_17_962 ();
 FILLCELL_X2 FILLER_0_17_1016 ();
 FILLCELL_X16 FILLER_0_17_1028 ();
 FILLCELL_X32 FILLER_0_17_1064 ();
 FILLCELL_X32 FILLER_0_17_1096 ();
 FILLCELL_X16 FILLER_0_17_1128 ();
 FILLCELL_X4 FILLER_0_17_1144 ();
 FILLCELL_X32 FILLER_0_18_1 ();
 FILLCELL_X32 FILLER_0_18_33 ();
 FILLCELL_X32 FILLER_0_18_65 ();
 FILLCELL_X32 FILLER_0_18_97 ();
 FILLCELL_X32 FILLER_0_18_129 ();
 FILLCELL_X32 FILLER_0_18_161 ();
 FILLCELL_X16 FILLER_0_18_193 ();
 FILLCELL_X8 FILLER_0_18_209 ();
 FILLCELL_X4 FILLER_0_18_217 ();
 FILLCELL_X2 FILLER_0_18_221 ();
 FILLCELL_X2 FILLER_0_18_298 ();
 FILLCELL_X1 FILLER_0_18_300 ();
 FILLCELL_X2 FILLER_0_18_341 ();
 FILLCELL_X2 FILLER_0_18_367 ();
 FILLCELL_X2 FILLER_0_18_376 ();
 FILLCELL_X4 FILLER_0_18_395 ();
 FILLCELL_X2 FILLER_0_18_402 ();
 FILLCELL_X1 FILLER_0_18_404 ();
 FILLCELL_X1 FILLER_0_18_409 ();
 FILLCELL_X1 FILLER_0_18_420 ();
 FILLCELL_X1 FILLER_0_18_448 ();
 FILLCELL_X2 FILLER_0_18_530 ();
 FILLCELL_X1 FILLER_0_18_549 ();
 FILLCELL_X2 FILLER_0_18_570 ();
 FILLCELL_X1 FILLER_0_18_572 ();
 FILLCELL_X1 FILLER_0_18_625 ();
 FILLCELL_X1 FILLER_0_18_639 ();
 FILLCELL_X1 FILLER_0_18_675 ();
 FILLCELL_X1 FILLER_0_18_686 ();
 FILLCELL_X1 FILLER_0_18_697 ();
 FILLCELL_X2 FILLER_0_18_708 ();
 FILLCELL_X2 FILLER_0_18_807 ();
 FILLCELL_X2 FILLER_0_18_822 ();
 FILLCELL_X1 FILLER_0_18_824 ();
 FILLCELL_X4 FILLER_0_18_829 ();
 FILLCELL_X2 FILLER_0_18_833 ();
 FILLCELL_X1 FILLER_0_18_835 ();
 FILLCELL_X2 FILLER_0_18_849 ();
 FILLCELL_X1 FILLER_0_18_851 ();
 FILLCELL_X8 FILLER_0_18_855 ();
 FILLCELL_X4 FILLER_0_18_863 ();
 FILLCELL_X2 FILLER_0_18_867 ();
 FILLCELL_X1 FILLER_0_18_869 ();
 FILLCELL_X2 FILLER_0_18_890 ();
 FILLCELL_X2 FILLER_0_18_903 ();
 FILLCELL_X2 FILLER_0_18_929 ();
 FILLCELL_X8 FILLER_0_18_956 ();
 FILLCELL_X4 FILLER_0_18_964 ();
 FILLCELL_X4 FILLER_0_18_978 ();
 FILLCELL_X1 FILLER_0_18_992 ();
 FILLCELL_X2 FILLER_0_18_998 ();
 FILLCELL_X2 FILLER_0_18_1020 ();
 FILLCELL_X1 FILLER_0_18_1031 ();
 FILLCELL_X1 FILLER_0_18_1042 ();
 FILLCELL_X32 FILLER_0_18_1058 ();
 FILLCELL_X32 FILLER_0_18_1090 ();
 FILLCELL_X16 FILLER_0_18_1122 ();
 FILLCELL_X8 FILLER_0_18_1138 ();
 FILLCELL_X2 FILLER_0_18_1146 ();
 FILLCELL_X32 FILLER_0_19_1 ();
 FILLCELL_X32 FILLER_0_19_33 ();
 FILLCELL_X32 FILLER_0_19_65 ();
 FILLCELL_X32 FILLER_0_19_97 ();
 FILLCELL_X32 FILLER_0_19_129 ();
 FILLCELL_X32 FILLER_0_19_161 ();
 FILLCELL_X16 FILLER_0_19_193 ();
 FILLCELL_X8 FILLER_0_19_209 ();
 FILLCELL_X1 FILLER_0_19_217 ();
 FILLCELL_X2 FILLER_0_19_254 ();
 FILLCELL_X1 FILLER_0_19_256 ();
 FILLCELL_X1 FILLER_0_19_267 ();
 FILLCELL_X4 FILLER_0_19_310 ();
 FILLCELL_X1 FILLER_0_19_335 ();
 FILLCELL_X2 FILLER_0_19_366 ();
 FILLCELL_X1 FILLER_0_19_381 ();
 FILLCELL_X1 FILLER_0_19_424 ();
 FILLCELL_X2 FILLER_0_19_456 ();
 FILLCELL_X2 FILLER_0_19_557 ();
 FILLCELL_X1 FILLER_0_19_559 ();
 FILLCELL_X1 FILLER_0_19_604 ();
 FILLCELL_X4 FILLER_0_19_639 ();
 FILLCELL_X1 FILLER_0_19_667 ();
 FILLCELL_X2 FILLER_0_19_678 ();
 FILLCELL_X1 FILLER_0_19_680 ();
 FILLCELL_X2 FILLER_0_19_704 ();
 FILLCELL_X1 FILLER_0_19_789 ();
 FILLCELL_X4 FILLER_0_19_800 ();
 FILLCELL_X2 FILLER_0_19_804 ();
 FILLCELL_X1 FILLER_0_19_806 ();
 FILLCELL_X2 FILLER_0_19_810 ();
 FILLCELL_X2 FILLER_0_19_830 ();
 FILLCELL_X1 FILLER_0_19_832 ();
 FILLCELL_X2 FILLER_0_19_857 ();
 FILLCELL_X4 FILLER_0_19_880 ();
 FILLCELL_X2 FILLER_0_19_884 ();
 FILLCELL_X2 FILLER_0_19_902 ();
 FILLCELL_X1 FILLER_0_19_904 ();
 FILLCELL_X8 FILLER_0_19_915 ();
 FILLCELL_X1 FILLER_0_19_962 ();
 FILLCELL_X2 FILLER_0_19_982 ();
 FILLCELL_X1 FILLER_0_19_984 ();
 FILLCELL_X8 FILLER_0_19_1005 ();
 FILLCELL_X1 FILLER_0_19_1013 ();
 FILLCELL_X32 FILLER_0_19_1049 ();
 FILLCELL_X32 FILLER_0_19_1081 ();
 FILLCELL_X32 FILLER_0_19_1113 ();
 FILLCELL_X2 FILLER_0_19_1145 ();
 FILLCELL_X1 FILLER_0_19_1147 ();
 FILLCELL_X32 FILLER_0_20_1 ();
 FILLCELL_X32 FILLER_0_20_33 ();
 FILLCELL_X32 FILLER_0_20_65 ();
 FILLCELL_X32 FILLER_0_20_97 ();
 FILLCELL_X32 FILLER_0_20_129 ();
 FILLCELL_X32 FILLER_0_20_161 ();
 FILLCELL_X16 FILLER_0_20_193 ();
 FILLCELL_X4 FILLER_0_20_209 ();
 FILLCELL_X2 FILLER_0_20_213 ();
 FILLCELL_X1 FILLER_0_20_240 ();
 FILLCELL_X2 FILLER_0_20_263 ();
 FILLCELL_X1 FILLER_0_20_265 ();
 FILLCELL_X2 FILLER_0_20_276 ();
 FILLCELL_X1 FILLER_0_20_278 ();
 FILLCELL_X1 FILLER_0_20_325 ();
 FILLCELL_X1 FILLER_0_20_346 ();
 FILLCELL_X4 FILLER_0_20_364 ();
 FILLCELL_X2 FILLER_0_20_368 ();
 FILLCELL_X1 FILLER_0_20_380 ();
 FILLCELL_X8 FILLER_0_20_391 ();
 FILLCELL_X4 FILLER_0_20_399 ();
 FILLCELL_X4 FILLER_0_20_406 ();
 FILLCELL_X1 FILLER_0_20_410 ();
 FILLCELL_X1 FILLER_0_20_414 ();
 FILLCELL_X2 FILLER_0_20_459 ();
 FILLCELL_X1 FILLER_0_20_500 ();
 FILLCELL_X2 FILLER_0_20_518 ();
 FILLCELL_X1 FILLER_0_20_545 ();
 FILLCELL_X1 FILLER_0_20_551 ();
 FILLCELL_X1 FILLER_0_20_558 ();
 FILLCELL_X1 FILLER_0_20_607 ();
 FILLCELL_X2 FILLER_0_20_625 ();
 FILLCELL_X1 FILLER_0_20_630 ();
 FILLCELL_X16 FILLER_0_20_632 ();
 FILLCELL_X8 FILLER_0_20_648 ();
 FILLCELL_X2 FILLER_0_20_685 ();
 FILLCELL_X1 FILLER_0_20_687 ();
 FILLCELL_X1 FILLER_0_20_703 ();
 FILLCELL_X2 FILLER_0_20_723 ();
 FILLCELL_X1 FILLER_0_20_725 ();
 FILLCELL_X1 FILLER_0_20_750 ();
 FILLCELL_X4 FILLER_0_20_763 ();
 FILLCELL_X1 FILLER_0_20_767 ();
 FILLCELL_X2 FILLER_0_20_778 ();
 FILLCELL_X1 FILLER_0_20_780 ();
 FILLCELL_X4 FILLER_0_20_788 ();
 FILLCELL_X1 FILLER_0_20_792 ();
 FILLCELL_X8 FILLER_0_20_797 ();
 FILLCELL_X2 FILLER_0_20_865 ();
 FILLCELL_X4 FILLER_0_20_881 ();
 FILLCELL_X4 FILLER_0_20_893 ();
 FILLCELL_X2 FILLER_0_20_897 ();
 FILLCELL_X8 FILLER_0_20_909 ();
 FILLCELL_X2 FILLER_0_20_917 ();
 FILLCELL_X1 FILLER_0_20_919 ();
 FILLCELL_X2 FILLER_0_20_993 ();
 FILLCELL_X1 FILLER_0_20_995 ();
 FILLCELL_X8 FILLER_0_20_1006 ();
 FILLCELL_X4 FILLER_0_20_1014 ();
 FILLCELL_X2 FILLER_0_20_1018 ();
 FILLCELL_X1 FILLER_0_20_1020 ();
 FILLCELL_X32 FILLER_0_20_1040 ();
 FILLCELL_X32 FILLER_0_20_1072 ();
 FILLCELL_X32 FILLER_0_20_1104 ();
 FILLCELL_X8 FILLER_0_20_1136 ();
 FILLCELL_X4 FILLER_0_20_1144 ();
 FILLCELL_X32 FILLER_0_21_1 ();
 FILLCELL_X32 FILLER_0_21_33 ();
 FILLCELL_X32 FILLER_0_21_65 ();
 FILLCELL_X32 FILLER_0_21_97 ();
 FILLCELL_X32 FILLER_0_21_129 ();
 FILLCELL_X32 FILLER_0_21_161 ();
 FILLCELL_X8 FILLER_0_21_193 ();
 FILLCELL_X4 FILLER_0_21_201 ();
 FILLCELL_X2 FILLER_0_21_220 ();
 FILLCELL_X8 FILLER_0_21_237 ();
 FILLCELL_X1 FILLER_0_21_245 ();
 FILLCELL_X2 FILLER_0_21_256 ();
 FILLCELL_X2 FILLER_0_21_268 ();
 FILLCELL_X2 FILLER_0_21_297 ();
 FILLCELL_X1 FILLER_0_21_299 ();
 FILLCELL_X4 FILLER_0_21_354 ();
 FILLCELL_X1 FILLER_0_21_358 ();
 FILLCELL_X8 FILLER_0_21_362 ();
 FILLCELL_X2 FILLER_0_21_370 ();
 FILLCELL_X1 FILLER_0_21_372 ();
 FILLCELL_X2 FILLER_0_21_375 ();
 FILLCELL_X2 FILLER_0_21_387 ();
 FILLCELL_X2 FILLER_0_21_418 ();
 FILLCELL_X1 FILLER_0_21_430 ();
 FILLCELL_X1 FILLER_0_21_438 ();
 FILLCELL_X1 FILLER_0_21_442 ();
 FILLCELL_X2 FILLER_0_21_465 ();
 FILLCELL_X1 FILLER_0_21_502 ();
 FILLCELL_X1 FILLER_0_21_518 ();
 FILLCELL_X1 FILLER_0_21_524 ();
 FILLCELL_X2 FILLER_0_21_535 ();
 FILLCELL_X1 FILLER_0_21_537 ();
 FILLCELL_X2 FILLER_0_21_560 ();
 FILLCELL_X1 FILLER_0_21_572 ();
 FILLCELL_X4 FILLER_0_21_576 ();
 FILLCELL_X16 FILLER_0_21_593 ();
 FILLCELL_X4 FILLER_0_21_609 ();
 FILLCELL_X16 FILLER_0_21_615 ();
 FILLCELL_X4 FILLER_0_21_631 ();
 FILLCELL_X2 FILLER_0_21_635 ();
 FILLCELL_X1 FILLER_0_21_637 ();
 FILLCELL_X8 FILLER_0_21_648 ();
 FILLCELL_X2 FILLER_0_21_673 ();
 FILLCELL_X1 FILLER_0_21_675 ();
 FILLCELL_X4 FILLER_0_21_685 ();
 FILLCELL_X1 FILLER_0_21_730 ();
 FILLCELL_X1 FILLER_0_21_741 ();
 FILLCELL_X8 FILLER_0_21_757 ();
 FILLCELL_X2 FILLER_0_21_775 ();
 FILLCELL_X2 FILLER_0_21_800 ();
 FILLCELL_X1 FILLER_0_21_802 ();
 FILLCELL_X1 FILLER_0_21_812 ();
 FILLCELL_X1 FILLER_0_21_825 ();
 FILLCELL_X1 FILLER_0_21_843 ();
 FILLCELL_X1 FILLER_0_21_850 ();
 FILLCELL_X4 FILLER_0_21_861 ();
 FILLCELL_X2 FILLER_0_21_865 ();
 FILLCELL_X2 FILLER_0_21_891 ();
 FILLCELL_X1 FILLER_0_21_893 ();
 FILLCELL_X4 FILLER_0_21_901 ();
 FILLCELL_X2 FILLER_0_21_905 ();
 FILLCELL_X1 FILLER_0_21_907 ();
 FILLCELL_X1 FILLER_0_21_910 ();
 FILLCELL_X16 FILLER_0_21_921 ();
 FILLCELL_X2 FILLER_0_21_937 ();
 FILLCELL_X2 FILLER_0_21_949 ();
 FILLCELL_X1 FILLER_0_21_966 ();
 FILLCELL_X2 FILLER_0_21_977 ();
 FILLCELL_X2 FILLER_0_21_988 ();
 FILLCELL_X2 FILLER_0_21_995 ();
 FILLCELL_X1 FILLER_0_21_997 ();
 FILLCELL_X8 FILLER_0_21_1008 ();
 FILLCELL_X4 FILLER_0_21_1016 ();
 FILLCELL_X1 FILLER_0_21_1030 ();
 FILLCELL_X8 FILLER_0_21_1036 ();
 FILLCELL_X4 FILLER_0_21_1044 ();
 FILLCELL_X1 FILLER_0_21_1048 ();
 FILLCELL_X32 FILLER_0_21_1059 ();
 FILLCELL_X32 FILLER_0_21_1091 ();
 FILLCELL_X16 FILLER_0_21_1123 ();
 FILLCELL_X8 FILLER_0_21_1139 ();
 FILLCELL_X1 FILLER_0_21_1147 ();
 FILLCELL_X32 FILLER_0_22_1 ();
 FILLCELL_X32 FILLER_0_22_33 ();
 FILLCELL_X32 FILLER_0_22_65 ();
 FILLCELL_X32 FILLER_0_22_97 ();
 FILLCELL_X32 FILLER_0_22_129 ();
 FILLCELL_X32 FILLER_0_22_161 ();
 FILLCELL_X16 FILLER_0_22_193 ();
 FILLCELL_X4 FILLER_0_22_209 ();
 FILLCELL_X2 FILLER_0_22_223 ();
 FILLCELL_X4 FILLER_0_22_244 ();
 FILLCELL_X1 FILLER_0_22_248 ();
 FILLCELL_X4 FILLER_0_22_269 ();
 FILLCELL_X2 FILLER_0_22_273 ();
 FILLCELL_X1 FILLER_0_22_275 ();
 FILLCELL_X1 FILLER_0_22_297 ();
 FILLCELL_X2 FILLER_0_22_308 ();
 FILLCELL_X2 FILLER_0_22_326 ();
 FILLCELL_X4 FILLER_0_22_347 ();
 FILLCELL_X1 FILLER_0_22_377 ();
 FILLCELL_X1 FILLER_0_22_434 ();
 FILLCELL_X1 FILLER_0_22_452 ();
 FILLCELL_X16 FILLER_0_22_463 ();
 FILLCELL_X8 FILLER_0_22_479 ();
 FILLCELL_X1 FILLER_0_22_492 ();
 FILLCELL_X1 FILLER_0_22_500 ();
 FILLCELL_X1 FILLER_0_22_511 ();
 FILLCELL_X1 FILLER_0_22_522 ();
 FILLCELL_X2 FILLER_0_22_527 ();
 FILLCELL_X4 FILLER_0_22_549 ();
 FILLCELL_X2 FILLER_0_22_570 ();
 FILLCELL_X2 FILLER_0_22_593 ();
 FILLCELL_X4 FILLER_0_22_625 ();
 FILLCELL_X2 FILLER_0_22_629 ();
 FILLCELL_X1 FILLER_0_22_632 ();
 FILLCELL_X16 FILLER_0_22_643 ();
 FILLCELL_X2 FILLER_0_22_684 ();
 FILLCELL_X1 FILLER_0_22_686 ();
 FILLCELL_X4 FILLER_0_22_697 ();
 FILLCELL_X2 FILLER_0_22_716 ();
 FILLCELL_X2 FILLER_0_22_733 ();
 FILLCELL_X1 FILLER_0_22_735 ();
 FILLCELL_X1 FILLER_0_22_746 ();
 FILLCELL_X8 FILLER_0_22_752 ();
 FILLCELL_X1 FILLER_0_22_797 ();
 FILLCELL_X2 FILLER_0_22_808 ();
 FILLCELL_X2 FILLER_0_22_840 ();
 FILLCELL_X1 FILLER_0_22_880 ();
 FILLCELL_X1 FILLER_0_22_891 ();
 FILLCELL_X1 FILLER_0_22_896 ();
 FILLCELL_X1 FILLER_0_22_907 ();
 FILLCELL_X16 FILLER_0_22_918 ();
 FILLCELL_X8 FILLER_0_22_934 ();
 FILLCELL_X4 FILLER_0_22_961 ();
 FILLCELL_X4 FILLER_0_22_985 ();
 FILLCELL_X4 FILLER_0_22_999 ();
 FILLCELL_X1 FILLER_0_22_1003 ();
 FILLCELL_X8 FILLER_0_22_1014 ();
 FILLCELL_X4 FILLER_0_22_1022 ();
 FILLCELL_X1 FILLER_0_22_1026 ();
 FILLCELL_X32 FILLER_0_22_1067 ();
 FILLCELL_X32 FILLER_0_22_1099 ();
 FILLCELL_X16 FILLER_0_22_1131 ();
 FILLCELL_X1 FILLER_0_22_1147 ();
 FILLCELL_X32 FILLER_0_23_1 ();
 FILLCELL_X32 FILLER_0_23_33 ();
 FILLCELL_X32 FILLER_0_23_65 ();
 FILLCELL_X32 FILLER_0_23_97 ();
 FILLCELL_X32 FILLER_0_23_129 ();
 FILLCELL_X32 FILLER_0_23_161 ();
 FILLCELL_X8 FILLER_0_23_193 ();
 FILLCELL_X4 FILLER_0_23_201 ();
 FILLCELL_X1 FILLER_0_23_205 ();
 FILLCELL_X2 FILLER_0_23_215 ();
 FILLCELL_X1 FILLER_0_23_217 ();
 FILLCELL_X1 FILLER_0_23_223 ();
 FILLCELL_X4 FILLER_0_23_234 ();
 FILLCELL_X2 FILLER_0_23_238 ();
 FILLCELL_X1 FILLER_0_23_240 ();
 FILLCELL_X8 FILLER_0_23_246 ();
 FILLCELL_X4 FILLER_0_23_254 ();
 FILLCELL_X1 FILLER_0_23_258 ();
 FILLCELL_X4 FILLER_0_23_264 ();
 FILLCELL_X1 FILLER_0_23_268 ();
 FILLCELL_X1 FILLER_0_23_279 ();
 FILLCELL_X1 FILLER_0_23_404 ();
 FILLCELL_X1 FILLER_0_23_415 ();
 FILLCELL_X2 FILLER_0_23_427 ();
 FILLCELL_X1 FILLER_0_23_460 ();
 FILLCELL_X2 FILLER_0_23_496 ();
 FILLCELL_X4 FILLER_0_23_512 ();
 FILLCELL_X1 FILLER_0_23_528 ();
 FILLCELL_X2 FILLER_0_23_539 ();
 FILLCELL_X2 FILLER_0_23_571 ();
 FILLCELL_X1 FILLER_0_23_573 ();
 FILLCELL_X1 FILLER_0_23_612 ();
 FILLCELL_X4 FILLER_0_23_632 ();
 FILLCELL_X2 FILLER_0_23_636 ();
 FILLCELL_X4 FILLER_0_23_660 ();
 FILLCELL_X2 FILLER_0_23_664 ();
 FILLCELL_X1 FILLER_0_23_678 ();
 FILLCELL_X16 FILLER_0_23_723 ();
 FILLCELL_X4 FILLER_0_23_739 ();
 FILLCELL_X2 FILLER_0_23_743 ();
 FILLCELL_X1 FILLER_0_23_745 ();
 FILLCELL_X1 FILLER_0_23_756 ();
 FILLCELL_X1 FILLER_0_23_798 ();
 FILLCELL_X2 FILLER_0_23_906 ();
 FILLCELL_X4 FILLER_0_23_913 ();
 FILLCELL_X1 FILLER_0_23_917 ();
 FILLCELL_X8 FILLER_0_23_928 ();
 FILLCELL_X2 FILLER_0_23_936 ();
 FILLCELL_X2 FILLER_0_23_975 ();
 FILLCELL_X2 FILLER_0_23_991 ();
 FILLCELL_X1 FILLER_0_23_993 ();
 FILLCELL_X8 FILLER_0_23_1004 ();
 FILLCELL_X2 FILLER_0_23_1012 ();
 FILLCELL_X2 FILLER_0_23_1029 ();
 FILLCELL_X2 FILLER_0_23_1046 ();
 FILLCELL_X32 FILLER_0_23_1078 ();
 FILLCELL_X32 FILLER_0_23_1110 ();
 FILLCELL_X4 FILLER_0_23_1142 ();
 FILLCELL_X2 FILLER_0_23_1146 ();
 FILLCELL_X32 FILLER_0_24_1 ();
 FILLCELL_X32 FILLER_0_24_33 ();
 FILLCELL_X32 FILLER_0_24_65 ();
 FILLCELL_X32 FILLER_0_24_97 ();
 FILLCELL_X32 FILLER_0_24_129 ();
 FILLCELL_X32 FILLER_0_24_161 ();
 FILLCELL_X8 FILLER_0_24_193 ();
 FILLCELL_X1 FILLER_0_24_201 ();
 FILLCELL_X4 FILLER_0_24_212 ();
 FILLCELL_X2 FILLER_0_24_254 ();
 FILLCELL_X2 FILLER_0_24_261 ();
 FILLCELL_X1 FILLER_0_24_263 ();
 FILLCELL_X1 FILLER_0_24_277 ();
 FILLCELL_X2 FILLER_0_24_298 ();
 FILLCELL_X1 FILLER_0_24_346 ();
 FILLCELL_X1 FILLER_0_24_381 ();
 FILLCELL_X8 FILLER_0_24_411 ();
 FILLCELL_X2 FILLER_0_24_429 ();
 FILLCELL_X2 FILLER_0_24_438 ();
 FILLCELL_X1 FILLER_0_24_447 ();
 FILLCELL_X1 FILLER_0_24_452 ();
 FILLCELL_X1 FILLER_0_24_467 ();
 FILLCELL_X1 FILLER_0_24_484 ();
 FILLCELL_X4 FILLER_0_24_502 ();
 FILLCELL_X1 FILLER_0_24_506 ();
 FILLCELL_X4 FILLER_0_24_517 ();
 FILLCELL_X2 FILLER_0_24_549 ();
 FILLCELL_X1 FILLER_0_24_551 ();
 FILLCELL_X8 FILLER_0_24_562 ();
 FILLCELL_X1 FILLER_0_24_570 ();
 FILLCELL_X4 FILLER_0_24_626 ();
 FILLCELL_X1 FILLER_0_24_630 ();
 FILLCELL_X8 FILLER_0_24_632 ();
 FILLCELL_X1 FILLER_0_24_663 ();
 FILLCELL_X2 FILLER_0_24_667 ();
 FILLCELL_X4 FILLER_0_24_685 ();
 FILLCELL_X8 FILLER_0_24_714 ();
 FILLCELL_X4 FILLER_0_24_742 ();
 FILLCELL_X1 FILLER_0_24_746 ();
 FILLCELL_X2 FILLER_0_24_765 ();
 FILLCELL_X2 FILLER_0_24_820 ();
 FILLCELL_X1 FILLER_0_24_828 ();
 FILLCELL_X1 FILLER_0_24_867 ();
 FILLCELL_X8 FILLER_0_24_899 ();
 FILLCELL_X2 FILLER_0_24_907 ();
 FILLCELL_X1 FILLER_0_24_909 ();
 FILLCELL_X2 FILLER_0_24_917 ();
 FILLCELL_X1 FILLER_0_24_924 ();
 FILLCELL_X2 FILLER_0_24_940 ();
 FILLCELL_X2 FILLER_0_24_957 ();
 FILLCELL_X1 FILLER_0_24_959 ();
 FILLCELL_X1 FILLER_0_24_965 ();
 FILLCELL_X4 FILLER_0_24_981 ();
 FILLCELL_X1 FILLER_0_24_1014 ();
 FILLCELL_X1 FILLER_0_24_1030 ();
 FILLCELL_X2 FILLER_0_24_1055 ();
 FILLCELL_X1 FILLER_0_24_1057 ();
 FILLCELL_X2 FILLER_0_24_1063 ();
 FILLCELL_X1 FILLER_0_24_1065 ();
 FILLCELL_X32 FILLER_0_24_1076 ();
 FILLCELL_X32 FILLER_0_24_1108 ();
 FILLCELL_X8 FILLER_0_24_1140 ();
 FILLCELL_X32 FILLER_0_25_1 ();
 FILLCELL_X32 FILLER_0_25_33 ();
 FILLCELL_X32 FILLER_0_25_65 ();
 FILLCELL_X32 FILLER_0_25_97 ();
 FILLCELL_X32 FILLER_0_25_129 ();
 FILLCELL_X32 FILLER_0_25_161 ();
 FILLCELL_X8 FILLER_0_25_193 ();
 FILLCELL_X4 FILLER_0_25_201 ();
 FILLCELL_X2 FILLER_0_25_205 ();
 FILLCELL_X1 FILLER_0_25_207 ();
 FILLCELL_X8 FILLER_0_25_218 ();
 FILLCELL_X2 FILLER_0_25_226 ();
 FILLCELL_X1 FILLER_0_25_228 ();
 FILLCELL_X2 FILLER_0_25_239 ();
 FILLCELL_X2 FILLER_0_25_271 ();
 FILLCELL_X1 FILLER_0_25_273 ();
 FILLCELL_X2 FILLER_0_25_284 ();
 FILLCELL_X1 FILLER_0_25_286 ();
 FILLCELL_X4 FILLER_0_25_292 ();
 FILLCELL_X2 FILLER_0_25_305 ();
 FILLCELL_X2 FILLER_0_25_317 ();
 FILLCELL_X1 FILLER_0_25_319 ();
 FILLCELL_X2 FILLER_0_25_362 ();
 FILLCELL_X1 FILLER_0_25_374 ();
 FILLCELL_X8 FILLER_0_25_399 ();
 FILLCELL_X1 FILLER_0_25_407 ();
 FILLCELL_X4 FILLER_0_25_418 ();
 FILLCELL_X2 FILLER_0_25_422 ();
 FILLCELL_X1 FILLER_0_25_443 ();
 FILLCELL_X1 FILLER_0_25_499 ();
 FILLCELL_X2 FILLER_0_25_510 ();
 FILLCELL_X1 FILLER_0_25_512 ();
 FILLCELL_X2 FILLER_0_25_545 ();
 FILLCELL_X4 FILLER_0_25_556 ();
 FILLCELL_X2 FILLER_0_25_560 ();
 FILLCELL_X1 FILLER_0_25_566 ();
 FILLCELL_X1 FILLER_0_25_569 ();
 FILLCELL_X2 FILLER_0_25_602 ();
 FILLCELL_X8 FILLER_0_25_628 ();
 FILLCELL_X4 FILLER_0_25_636 ();
 FILLCELL_X2 FILLER_0_25_640 ();
 FILLCELL_X1 FILLER_0_25_652 ();
 FILLCELL_X4 FILLER_0_25_659 ();
 FILLCELL_X16 FILLER_0_25_673 ();
 FILLCELL_X1 FILLER_0_25_689 ();
 FILLCELL_X2 FILLER_0_25_699 ();
 FILLCELL_X1 FILLER_0_25_701 ();
 FILLCELL_X2 FILLER_0_25_719 ();
 FILLCELL_X1 FILLER_0_25_727 ();
 FILLCELL_X1 FILLER_0_25_738 ();
 FILLCELL_X1 FILLER_0_25_749 ();
 FILLCELL_X1 FILLER_0_25_755 ();
 FILLCELL_X1 FILLER_0_25_766 ();
 FILLCELL_X8 FILLER_0_25_791 ();
 FILLCELL_X2 FILLER_0_25_799 ();
 FILLCELL_X1 FILLER_0_25_801 ();
 FILLCELL_X1 FILLER_0_25_874 ();
 FILLCELL_X1 FILLER_0_25_882 ();
 FILLCELL_X1 FILLER_0_25_935 ();
 FILLCELL_X1 FILLER_0_25_998 ();
 FILLCELL_X2 FILLER_0_25_1030 ();
 FILLCELL_X2 FILLER_0_25_1037 ();
 FILLCELL_X1 FILLER_0_25_1039 ();
 FILLCELL_X1 FILLER_0_25_1069 ();
 FILLCELL_X2 FILLER_0_25_1079 ();
 FILLCELL_X32 FILLER_0_25_1091 ();
 FILLCELL_X16 FILLER_0_25_1123 ();
 FILLCELL_X8 FILLER_0_25_1139 ();
 FILLCELL_X1 FILLER_0_25_1147 ();
 FILLCELL_X32 FILLER_0_26_1 ();
 FILLCELL_X32 FILLER_0_26_33 ();
 FILLCELL_X32 FILLER_0_26_65 ();
 FILLCELL_X32 FILLER_0_26_97 ();
 FILLCELL_X32 FILLER_0_26_129 ();
 FILLCELL_X32 FILLER_0_26_161 ();
 FILLCELL_X4 FILLER_0_26_193 ();
 FILLCELL_X1 FILLER_0_26_197 ();
 FILLCELL_X32 FILLER_0_26_203 ();
 FILLCELL_X1 FILLER_0_26_255 ();
 FILLCELL_X4 FILLER_0_26_261 ();
 FILLCELL_X2 FILLER_0_26_270 ();
 FILLCELL_X2 FILLER_0_26_282 ();
 FILLCELL_X1 FILLER_0_26_284 ();
 FILLCELL_X2 FILLER_0_26_295 ();
 FILLCELL_X1 FILLER_0_26_297 ();
 FILLCELL_X2 FILLER_0_26_308 ();
 FILLCELL_X1 FILLER_0_26_310 ();
 FILLCELL_X4 FILLER_0_26_321 ();
 FILLCELL_X2 FILLER_0_26_338 ();
 FILLCELL_X1 FILLER_0_26_340 ();
 FILLCELL_X2 FILLER_0_26_367 ();
 FILLCELL_X1 FILLER_0_26_402 ();
 FILLCELL_X1 FILLER_0_26_467 ();
 FILLCELL_X2 FILLER_0_26_526 ();
 FILLCELL_X1 FILLER_0_26_528 ();
 FILLCELL_X2 FILLER_0_26_556 ();
 FILLCELL_X2 FILLER_0_26_589 ();
 FILLCELL_X2 FILLER_0_26_601 ();
 FILLCELL_X1 FILLER_0_26_603 ();
 FILLCELL_X1 FILLER_0_26_630 ();
 FILLCELL_X1 FILLER_0_26_671 ();
 FILLCELL_X8 FILLER_0_26_699 ();
 FILLCELL_X2 FILLER_0_26_707 ();
 FILLCELL_X1 FILLER_0_26_709 ();
 FILLCELL_X4 FILLER_0_26_720 ();
 FILLCELL_X2 FILLER_0_26_724 ();
 FILLCELL_X8 FILLER_0_26_761 ();
 FILLCELL_X1 FILLER_0_26_769 ();
 FILLCELL_X2 FILLER_0_26_777 ();
 FILLCELL_X1 FILLER_0_26_786 ();
 FILLCELL_X2 FILLER_0_26_794 ();
 FILLCELL_X1 FILLER_0_26_800 ();
 FILLCELL_X1 FILLER_0_26_811 ();
 FILLCELL_X4 FILLER_0_26_854 ();
 FILLCELL_X1 FILLER_0_26_858 ();
 FILLCELL_X4 FILLER_0_26_862 ();
 FILLCELL_X1 FILLER_0_26_866 ();
 FILLCELL_X2 FILLER_0_26_931 ();
 FILLCELL_X4 FILLER_0_26_943 ();
 FILLCELL_X1 FILLER_0_26_954 ();
 FILLCELL_X2 FILLER_0_26_965 ();
 FILLCELL_X1 FILLER_0_26_967 ();
 FILLCELL_X2 FILLER_0_26_978 ();
 FILLCELL_X2 FILLER_0_26_1011 ();
 FILLCELL_X1 FILLER_0_26_1028 ();
 FILLCELL_X4 FILLER_0_26_1059 ();
 FILLCELL_X2 FILLER_0_26_1068 ();
 FILLCELL_X32 FILLER_0_26_1080 ();
 FILLCELL_X32 FILLER_0_26_1112 ();
 FILLCELL_X4 FILLER_0_26_1144 ();
 FILLCELL_X32 FILLER_0_27_1 ();
 FILLCELL_X32 FILLER_0_27_33 ();
 FILLCELL_X32 FILLER_0_27_65 ();
 FILLCELL_X32 FILLER_0_27_97 ();
 FILLCELL_X32 FILLER_0_27_129 ();
 FILLCELL_X32 FILLER_0_27_161 ();
 FILLCELL_X2 FILLER_0_27_193 ();
 FILLCELL_X4 FILLER_0_27_205 ();
 FILLCELL_X1 FILLER_0_27_229 ();
 FILLCELL_X8 FILLER_0_27_272 ();
 FILLCELL_X4 FILLER_0_27_280 ();
 FILLCELL_X8 FILLER_0_27_308 ();
 FILLCELL_X2 FILLER_0_27_316 ();
 FILLCELL_X1 FILLER_0_27_318 ();
 FILLCELL_X4 FILLER_0_27_347 ();
 FILLCELL_X2 FILLER_0_27_364 ();
 FILLCELL_X2 FILLER_0_27_379 ();
 FILLCELL_X2 FILLER_0_27_418 ();
 FILLCELL_X1 FILLER_0_27_420 ();
 FILLCELL_X1 FILLER_0_27_434 ();
 FILLCELL_X1 FILLER_0_27_526 ();
 FILLCELL_X1 FILLER_0_27_550 ();
 FILLCELL_X2 FILLER_0_27_592 ();
 FILLCELL_X4 FILLER_0_27_606 ();
 FILLCELL_X1 FILLER_0_27_619 ();
 FILLCELL_X8 FILLER_0_27_668 ();
 FILLCELL_X2 FILLER_0_27_692 ();
 FILLCELL_X1 FILLER_0_27_694 ();
 FILLCELL_X2 FILLER_0_27_712 ();
 FILLCELL_X1 FILLER_0_27_714 ();
 FILLCELL_X2 FILLER_0_27_758 ();
 FILLCELL_X1 FILLER_0_27_760 ();
 FILLCELL_X4 FILLER_0_27_775 ();
 FILLCELL_X2 FILLER_0_27_779 ();
 FILLCELL_X4 FILLER_0_27_795 ();
 FILLCELL_X1 FILLER_0_27_799 ();
 FILLCELL_X1 FILLER_0_27_813 ();
 FILLCELL_X2 FILLER_0_27_827 ();
 FILLCELL_X2 FILLER_0_27_873 ();
 FILLCELL_X1 FILLER_0_27_885 ();
 FILLCELL_X1 FILLER_0_27_890 ();
 FILLCELL_X1 FILLER_0_27_906 ();
 FILLCELL_X2 FILLER_0_27_931 ();
 FILLCELL_X1 FILLER_0_27_955 ();
 FILLCELL_X2 FILLER_0_27_966 ();
 FILLCELL_X2 FILLER_0_27_978 ();
 FILLCELL_X1 FILLER_0_27_980 ();
 FILLCELL_X1 FILLER_0_27_991 ();
 FILLCELL_X2 FILLER_0_27_1002 ();
 FILLCELL_X1 FILLER_0_27_1004 ();
 FILLCELL_X1 FILLER_0_27_1025 ();
 FILLCELL_X2 FILLER_0_27_1061 ();
 FILLCELL_X32 FILLER_0_27_1073 ();
 FILLCELL_X32 FILLER_0_27_1105 ();
 FILLCELL_X8 FILLER_0_27_1137 ();
 FILLCELL_X2 FILLER_0_27_1145 ();
 FILLCELL_X1 FILLER_0_27_1147 ();
 FILLCELL_X32 FILLER_0_28_1 ();
 FILLCELL_X32 FILLER_0_28_33 ();
 FILLCELL_X32 FILLER_0_28_65 ();
 FILLCELL_X32 FILLER_0_28_97 ();
 FILLCELL_X32 FILLER_0_28_129 ();
 FILLCELL_X32 FILLER_0_28_161 ();
 FILLCELL_X4 FILLER_0_28_193 ();
 FILLCELL_X4 FILLER_0_28_227 ();
 FILLCELL_X1 FILLER_0_28_256 ();
 FILLCELL_X2 FILLER_0_28_267 ();
 FILLCELL_X1 FILLER_0_28_269 ();
 FILLCELL_X2 FILLER_0_28_305 ();
 FILLCELL_X1 FILLER_0_28_317 ();
 FILLCELL_X1 FILLER_0_28_322 ();
 FILLCELL_X2 FILLER_0_28_357 ();
 FILLCELL_X4 FILLER_0_28_372 ();
 FILLCELL_X1 FILLER_0_28_441 ();
 FILLCELL_X2 FILLER_0_28_579 ();
 FILLCELL_X1 FILLER_0_28_586 ();
 FILLCELL_X2 FILLER_0_28_701 ();
 FILLCELL_X1 FILLER_0_28_703 ();
 FILLCELL_X4 FILLER_0_28_708 ();
 FILLCELL_X4 FILLER_0_28_725 ();
 FILLCELL_X1 FILLER_0_28_729 ();
 FILLCELL_X2 FILLER_0_28_768 ();
 FILLCELL_X1 FILLER_0_28_770 ();
 FILLCELL_X2 FILLER_0_28_774 ();
 FILLCELL_X2 FILLER_0_28_780 ();
 FILLCELL_X1 FILLER_0_28_782 ();
 FILLCELL_X4 FILLER_0_28_796 ();
 FILLCELL_X2 FILLER_0_28_800 ();
 FILLCELL_X2 FILLER_0_28_832 ();
 FILLCELL_X1 FILLER_0_28_858 ();
 FILLCELL_X4 FILLER_0_28_941 ();
 FILLCELL_X2 FILLER_0_28_990 ();
 FILLCELL_X1 FILLER_0_28_992 ();
 FILLCELL_X4 FILLER_0_28_1018 ();
 FILLCELL_X2 FILLER_0_28_1039 ();
 FILLCELL_X1 FILLER_0_28_1041 ();
 FILLCELL_X32 FILLER_0_28_1081 ();
 FILLCELL_X32 FILLER_0_28_1113 ();
 FILLCELL_X2 FILLER_0_28_1145 ();
 FILLCELL_X1 FILLER_0_28_1147 ();
 FILLCELL_X32 FILLER_0_29_1 ();
 FILLCELL_X32 FILLER_0_29_33 ();
 FILLCELL_X32 FILLER_0_29_65 ();
 FILLCELL_X32 FILLER_0_29_97 ();
 FILLCELL_X32 FILLER_0_29_129 ();
 FILLCELL_X16 FILLER_0_29_161 ();
 FILLCELL_X4 FILLER_0_29_177 ();
 FILLCELL_X2 FILLER_0_29_211 ();
 FILLCELL_X1 FILLER_0_29_242 ();
 FILLCELL_X1 FILLER_0_29_268 ();
 FILLCELL_X2 FILLER_0_29_279 ();
 FILLCELL_X2 FILLER_0_29_325 ();
 FILLCELL_X1 FILLER_0_29_327 ();
 FILLCELL_X1 FILLER_0_29_361 ();
 FILLCELL_X8 FILLER_0_29_371 ();
 FILLCELL_X2 FILLER_0_29_379 ();
 FILLCELL_X1 FILLER_0_29_381 ();
 FILLCELL_X1 FILLER_0_29_459 ();
 FILLCELL_X1 FILLER_0_29_499 ();
 FILLCELL_X1 FILLER_0_29_547 ();
 FILLCELL_X1 FILLER_0_29_607 ();
 FILLCELL_X2 FILLER_0_29_655 ();
 FILLCELL_X2 FILLER_0_29_671 ();
 FILLCELL_X1 FILLER_0_29_703 ();
 FILLCELL_X1 FILLER_0_29_718 ();
 FILLCELL_X2 FILLER_0_29_724 ();
 FILLCELL_X1 FILLER_0_29_726 ();
 FILLCELL_X8 FILLER_0_29_760 ();
 FILLCELL_X4 FILLER_0_29_768 ();
 FILLCELL_X16 FILLER_0_29_782 ();
 FILLCELL_X4 FILLER_0_29_798 ();
 FILLCELL_X1 FILLER_0_29_802 ();
 FILLCELL_X2 FILLER_0_29_834 ();
 FILLCELL_X8 FILLER_0_29_843 ();
 FILLCELL_X4 FILLER_0_29_851 ();
 FILLCELL_X2 FILLER_0_29_855 ();
 FILLCELL_X1 FILLER_0_29_857 ();
 FILLCELL_X1 FILLER_0_29_862 ();
 FILLCELL_X2 FILLER_0_29_887 ();
 FILLCELL_X2 FILLER_0_29_918 ();
 FILLCELL_X1 FILLER_0_29_969 ();
 FILLCELL_X1 FILLER_0_29_1020 ();
 FILLCELL_X2 FILLER_0_29_1033 ();
 FILLCELL_X1 FILLER_0_29_1054 ();
 FILLCELL_X2 FILLER_0_29_1080 ();
 FILLCELL_X1 FILLER_0_29_1082 ();
 FILLCELL_X32 FILLER_0_29_1093 ();
 FILLCELL_X16 FILLER_0_29_1125 ();
 FILLCELL_X4 FILLER_0_29_1141 ();
 FILLCELL_X2 FILLER_0_29_1145 ();
 FILLCELL_X1 FILLER_0_29_1147 ();
 FILLCELL_X32 FILLER_0_30_1 ();
 FILLCELL_X32 FILLER_0_30_33 ();
 FILLCELL_X32 FILLER_0_30_65 ();
 FILLCELL_X32 FILLER_0_30_97 ();
 FILLCELL_X32 FILLER_0_30_129 ();
 FILLCELL_X16 FILLER_0_30_161 ();
 FILLCELL_X1 FILLER_0_30_177 ();
 FILLCELL_X4 FILLER_0_30_198 ();
 FILLCELL_X1 FILLER_0_30_202 ();
 FILLCELL_X1 FILLER_0_30_223 ();
 FILLCELL_X1 FILLER_0_30_255 ();
 FILLCELL_X2 FILLER_0_30_271 ();
 FILLCELL_X1 FILLER_0_30_309 ();
 FILLCELL_X2 FILLER_0_30_333 ();
 FILLCELL_X1 FILLER_0_30_335 ();
 FILLCELL_X8 FILLER_0_30_339 ();
 FILLCELL_X2 FILLER_0_30_347 ();
 FILLCELL_X1 FILLER_0_30_365 ();
 FILLCELL_X16 FILLER_0_30_373 ();
 FILLCELL_X2 FILLER_0_30_389 ();
 FILLCELL_X1 FILLER_0_30_391 ();
 FILLCELL_X1 FILLER_0_30_435 ();
 FILLCELL_X1 FILLER_0_30_514 ();
 FILLCELL_X2 FILLER_0_30_568 ();
 FILLCELL_X1 FILLER_0_30_639 ();
 FILLCELL_X1 FILLER_0_30_664 ();
 FILLCELL_X1 FILLER_0_30_681 ();
 FILLCELL_X1 FILLER_0_30_692 ();
 FILLCELL_X2 FILLER_0_30_713 ();
 FILLCELL_X2 FILLER_0_30_737 ();
 FILLCELL_X1 FILLER_0_30_739 ();
 FILLCELL_X4 FILLER_0_30_747 ();
 FILLCELL_X4 FILLER_0_30_761 ();
 FILLCELL_X8 FILLER_0_30_769 ();
 FILLCELL_X4 FILLER_0_30_777 ();
 FILLCELL_X1 FILLER_0_30_781 ();
 FILLCELL_X4 FILLER_0_30_785 ();
 FILLCELL_X1 FILLER_0_30_789 ();
 FILLCELL_X2 FILLER_0_30_794 ();
 FILLCELL_X1 FILLER_0_30_805 ();
 FILLCELL_X8 FILLER_0_30_844 ();
 FILLCELL_X2 FILLER_0_30_852 ();
 FILLCELL_X2 FILLER_0_30_869 ();
 FILLCELL_X4 FILLER_0_30_946 ();
 FILLCELL_X1 FILLER_0_30_984 ();
 FILLCELL_X2 FILLER_0_30_995 ();
 FILLCELL_X1 FILLER_0_30_997 ();
 FILLCELL_X4 FILLER_0_30_1079 ();
 FILLCELL_X32 FILLER_0_30_1093 ();
 FILLCELL_X16 FILLER_0_30_1125 ();
 FILLCELL_X4 FILLER_0_30_1141 ();
 FILLCELL_X2 FILLER_0_30_1145 ();
 FILLCELL_X1 FILLER_0_30_1147 ();
 FILLCELL_X32 FILLER_0_31_1 ();
 FILLCELL_X32 FILLER_0_31_33 ();
 FILLCELL_X32 FILLER_0_31_65 ();
 FILLCELL_X32 FILLER_0_31_97 ();
 FILLCELL_X32 FILLER_0_31_129 ();
 FILLCELL_X8 FILLER_0_31_161 ();
 FILLCELL_X4 FILLER_0_31_179 ();
 FILLCELL_X2 FILLER_0_31_226 ();
 FILLCELL_X1 FILLER_0_31_228 ();
 FILLCELL_X2 FILLER_0_31_246 ();
 FILLCELL_X1 FILLER_0_31_248 ();
 FILLCELL_X1 FILLER_0_31_280 ();
 FILLCELL_X1 FILLER_0_31_307 ();
 FILLCELL_X2 FILLER_0_31_318 ();
 FILLCELL_X1 FILLER_0_31_320 ();
 FILLCELL_X2 FILLER_0_31_342 ();
 FILLCELL_X2 FILLER_0_31_355 ();
 FILLCELL_X8 FILLER_0_31_389 ();
 FILLCELL_X2 FILLER_0_31_397 ();
 FILLCELL_X2 FILLER_0_31_420 ();
 FILLCELL_X2 FILLER_0_31_640 ();
 FILLCELL_X1 FILLER_0_31_688 ();
 FILLCELL_X1 FILLER_0_31_696 ();
 FILLCELL_X1 FILLER_0_31_730 ();
 FILLCELL_X16 FILLER_0_31_747 ();
 FILLCELL_X1 FILLER_0_31_763 ();
 FILLCELL_X4 FILLER_0_31_778 ();
 FILLCELL_X1 FILLER_0_31_782 ();
 FILLCELL_X2 FILLER_0_31_834 ();
 FILLCELL_X1 FILLER_0_31_938 ();
 FILLCELL_X2 FILLER_0_31_949 ();
 FILLCELL_X1 FILLER_0_31_983 ();
 FILLCELL_X1 FILLER_0_31_1001 ();
 FILLCELL_X1 FILLER_0_31_1012 ();
 FILLCELL_X2 FILLER_0_31_1028 ();
 FILLCELL_X2 FILLER_0_31_1040 ();
 FILLCELL_X8 FILLER_0_31_1052 ();
 FILLCELL_X4 FILLER_0_31_1070 ();
 FILLCELL_X1 FILLER_0_31_1074 ();
 FILLCELL_X32 FILLER_0_31_1085 ();
 FILLCELL_X16 FILLER_0_31_1117 ();
 FILLCELL_X8 FILLER_0_31_1133 ();
 FILLCELL_X4 FILLER_0_31_1141 ();
 FILLCELL_X2 FILLER_0_31_1145 ();
 FILLCELL_X1 FILLER_0_31_1147 ();
 FILLCELL_X32 FILLER_0_32_1 ();
 FILLCELL_X32 FILLER_0_32_33 ();
 FILLCELL_X32 FILLER_0_32_65 ();
 FILLCELL_X32 FILLER_0_32_97 ();
 FILLCELL_X32 FILLER_0_32_129 ();
 FILLCELL_X8 FILLER_0_32_161 ();
 FILLCELL_X2 FILLER_0_32_169 ();
 FILLCELL_X1 FILLER_0_32_171 ();
 FILLCELL_X2 FILLER_0_32_182 ();
 FILLCELL_X1 FILLER_0_32_184 ();
 FILLCELL_X1 FILLER_0_32_190 ();
 FILLCELL_X4 FILLER_0_32_218 ();
 FILLCELL_X4 FILLER_0_32_232 ();
 FILLCELL_X4 FILLER_0_32_256 ();
 FILLCELL_X1 FILLER_0_32_277 ();
 FILLCELL_X2 FILLER_0_32_315 ();
 FILLCELL_X1 FILLER_0_32_347 ();
 FILLCELL_X1 FILLER_0_32_365 ();
 FILLCELL_X2 FILLER_0_32_383 ();
 FILLCELL_X1 FILLER_0_32_385 ();
 FILLCELL_X1 FILLER_0_32_409 ();
 FILLCELL_X1 FILLER_0_32_473 ();
 FILLCELL_X1 FILLER_0_32_503 ();
 FILLCELL_X1 FILLER_0_32_516 ();
 FILLCELL_X2 FILLER_0_32_639 ();
 FILLCELL_X1 FILLER_0_32_677 ();
 FILLCELL_X1 FILLER_0_32_693 ();
 FILLCELL_X1 FILLER_0_32_738 ();
 FILLCELL_X4 FILLER_0_32_755 ();
 FILLCELL_X2 FILLER_0_32_763 ();
 FILLCELL_X1 FILLER_0_32_765 ();
 FILLCELL_X1 FILLER_0_32_795 ();
 FILLCELL_X2 FILLER_0_32_834 ();
 FILLCELL_X4 FILLER_0_32_843 ();
 FILLCELL_X2 FILLER_0_32_847 ();
 FILLCELL_X1 FILLER_0_32_849 ();
 FILLCELL_X2 FILLER_0_32_865 ();
 FILLCELL_X1 FILLER_0_32_944 ();
 FILLCELL_X4 FILLER_0_32_955 ();
 FILLCELL_X1 FILLER_0_32_1000 ();
 FILLCELL_X8 FILLER_0_32_1052 ();
 FILLCELL_X1 FILLER_0_32_1060 ();
 FILLCELL_X32 FILLER_0_32_1071 ();
 FILLCELL_X32 FILLER_0_32_1103 ();
 FILLCELL_X8 FILLER_0_32_1135 ();
 FILLCELL_X4 FILLER_0_32_1143 ();
 FILLCELL_X1 FILLER_0_32_1147 ();
 FILLCELL_X32 FILLER_0_33_1 ();
 FILLCELL_X32 FILLER_0_33_33 ();
 FILLCELL_X32 FILLER_0_33_65 ();
 FILLCELL_X32 FILLER_0_33_97 ();
 FILLCELL_X16 FILLER_0_33_129 ();
 FILLCELL_X8 FILLER_0_33_145 ();
 FILLCELL_X4 FILLER_0_33_153 ();
 FILLCELL_X2 FILLER_0_33_157 ();
 FILLCELL_X1 FILLER_0_33_159 ();
 FILLCELL_X2 FILLER_0_33_175 ();
 FILLCELL_X2 FILLER_0_33_197 ();
 FILLCELL_X1 FILLER_0_33_199 ();
 FILLCELL_X2 FILLER_0_33_227 ();
 FILLCELL_X1 FILLER_0_33_229 ();
 FILLCELL_X2 FILLER_0_33_261 ();
 FILLCELL_X1 FILLER_0_33_263 ();
 FILLCELL_X2 FILLER_0_33_274 ();
 FILLCELL_X1 FILLER_0_33_276 ();
 FILLCELL_X2 FILLER_0_33_296 ();
 FILLCELL_X1 FILLER_0_33_298 ();
 FILLCELL_X1 FILLER_0_33_347 ();
 FILLCELL_X1 FILLER_0_33_389 ();
 FILLCELL_X4 FILLER_0_33_394 ();
 FILLCELL_X1 FILLER_0_33_398 ();
 FILLCELL_X1 FILLER_0_33_402 ();
 FILLCELL_X1 FILLER_0_33_456 ();
 FILLCELL_X1 FILLER_0_33_475 ();
 FILLCELL_X1 FILLER_0_33_537 ();
 FILLCELL_X1 FILLER_0_33_637 ();
 FILLCELL_X1 FILLER_0_33_663 ();
 FILLCELL_X1 FILLER_0_33_740 ();
 FILLCELL_X1 FILLER_0_33_748 ();
 FILLCELL_X4 FILLER_0_33_773 ();
 FILLCELL_X1 FILLER_0_33_777 ();
 FILLCELL_X2 FILLER_0_33_811 ();
 FILLCELL_X2 FILLER_0_33_840 ();
 FILLCELL_X1 FILLER_0_33_842 ();
 FILLCELL_X1 FILLER_0_33_853 ();
 FILLCELL_X1 FILLER_0_33_892 ();
 FILLCELL_X4 FILLER_0_33_959 ();
 FILLCELL_X2 FILLER_0_33_983 ();
 FILLCELL_X2 FILLER_0_33_1019 ();
 FILLCELL_X1 FILLER_0_33_1021 ();
 FILLCELL_X8 FILLER_0_33_1047 ();
 FILLCELL_X4 FILLER_0_33_1055 ();
 FILLCELL_X2 FILLER_0_33_1059 ();
 FILLCELL_X1 FILLER_0_33_1061 ();
 FILLCELL_X1 FILLER_0_33_1067 ();
 FILLCELL_X4 FILLER_0_33_1078 ();
 FILLCELL_X32 FILLER_0_33_1092 ();
 FILLCELL_X16 FILLER_0_33_1124 ();
 FILLCELL_X8 FILLER_0_33_1140 ();
 FILLCELL_X32 FILLER_0_34_1 ();
 FILLCELL_X32 FILLER_0_34_33 ();
 FILLCELL_X32 FILLER_0_34_65 ();
 FILLCELL_X32 FILLER_0_34_97 ();
 FILLCELL_X32 FILLER_0_34_129 ();
 FILLCELL_X8 FILLER_0_34_161 ();
 FILLCELL_X4 FILLER_0_34_169 ();
 FILLCELL_X2 FILLER_0_34_173 ();
 FILLCELL_X1 FILLER_0_34_217 ();
 FILLCELL_X2 FILLER_0_34_257 ();
 FILLCELL_X2 FILLER_0_34_310 ();
 FILLCELL_X1 FILLER_0_34_312 ();
 FILLCELL_X4 FILLER_0_34_384 ();
 FILLCELL_X1 FILLER_0_34_388 ();
 FILLCELL_X1 FILLER_0_34_399 ();
 FILLCELL_X1 FILLER_0_34_418 ();
 FILLCELL_X2 FILLER_0_34_433 ();
 FILLCELL_X1 FILLER_0_34_469 ();
 FILLCELL_X2 FILLER_0_34_664 ();
 FILLCELL_X2 FILLER_0_34_686 ();
 FILLCELL_X1 FILLER_0_34_688 ();
 FILLCELL_X2 FILLER_0_34_696 ();
 FILLCELL_X1 FILLER_0_34_698 ();
 FILLCELL_X8 FILLER_0_34_777 ();
 FILLCELL_X2 FILLER_0_34_785 ();
 FILLCELL_X2 FILLER_0_34_831 ();
 FILLCELL_X1 FILLER_0_34_833 ();
 FILLCELL_X1 FILLER_0_34_844 ();
 FILLCELL_X2 FILLER_0_34_858 ();
 FILLCELL_X2 FILLER_0_34_865 ();
 FILLCELL_X1 FILLER_0_34_867 ();
 FILLCELL_X2 FILLER_0_34_963 ();
 FILLCELL_X2 FILLER_0_34_975 ();
 FILLCELL_X1 FILLER_0_34_977 ();
 FILLCELL_X2 FILLER_0_34_985 ();
 FILLCELL_X2 FILLER_0_34_1011 ();
 FILLCELL_X2 FILLER_0_34_1028 ();
 FILLCELL_X8 FILLER_0_34_1053 ();
 FILLCELL_X1 FILLER_0_34_1061 ();
 FILLCELL_X2 FILLER_0_34_1077 ();
 FILLCELL_X1 FILLER_0_34_1079 ();
 FILLCELL_X32 FILLER_0_34_1090 ();
 FILLCELL_X16 FILLER_0_34_1122 ();
 FILLCELL_X8 FILLER_0_34_1138 ();
 FILLCELL_X2 FILLER_0_34_1146 ();
 FILLCELL_X32 FILLER_0_35_1 ();
 FILLCELL_X32 FILLER_0_35_33 ();
 FILLCELL_X32 FILLER_0_35_65 ();
 FILLCELL_X32 FILLER_0_35_97 ();
 FILLCELL_X16 FILLER_0_35_129 ();
 FILLCELL_X8 FILLER_0_35_145 ();
 FILLCELL_X4 FILLER_0_35_153 ();
 FILLCELL_X2 FILLER_0_35_157 ();
 FILLCELL_X1 FILLER_0_35_159 ();
 FILLCELL_X8 FILLER_0_35_165 ();
 FILLCELL_X4 FILLER_0_35_173 ();
 FILLCELL_X2 FILLER_0_35_177 ();
 FILLCELL_X2 FILLER_0_35_224 ();
 FILLCELL_X1 FILLER_0_35_226 ();
 FILLCELL_X1 FILLER_0_35_244 ();
 FILLCELL_X2 FILLER_0_35_281 ();
 FILLCELL_X1 FILLER_0_35_283 ();
 FILLCELL_X2 FILLER_0_35_291 ();
 FILLCELL_X1 FILLER_0_35_293 ();
 FILLCELL_X1 FILLER_0_35_304 ();
 FILLCELL_X1 FILLER_0_35_331 ();
 FILLCELL_X1 FILLER_0_35_339 ();
 FILLCELL_X16 FILLER_0_35_376 ();
 FILLCELL_X4 FILLER_0_35_392 ();
 FILLCELL_X1 FILLER_0_35_426 ();
 FILLCELL_X1 FILLER_0_35_470 ();
 FILLCELL_X2 FILLER_0_35_480 ();
 FILLCELL_X1 FILLER_0_35_661 ();
 FILLCELL_X2 FILLER_0_35_679 ();
 FILLCELL_X2 FILLER_0_35_706 ();
 FILLCELL_X1 FILLER_0_35_708 ();
 FILLCELL_X8 FILLER_0_35_769 ();
 FILLCELL_X4 FILLER_0_35_777 ();
 FILLCELL_X2 FILLER_0_35_781 ();
 FILLCELL_X2 FILLER_0_35_793 ();
 FILLCELL_X1 FILLER_0_35_808 ();
 FILLCELL_X2 FILLER_0_35_823 ();
 FILLCELL_X2 FILLER_0_35_840 ();
 FILLCELL_X2 FILLER_0_35_892 ();
 FILLCELL_X1 FILLER_0_35_909 ();
 FILLCELL_X1 FILLER_0_35_920 ();
 FILLCELL_X1 FILLER_0_35_945 ();
 FILLCELL_X2 FILLER_0_35_980 ();
 FILLCELL_X1 FILLER_0_35_1009 ();
 FILLCELL_X1 FILLER_0_35_1020 ();
 FILLCELL_X4 FILLER_0_35_1051 ();
 FILLCELL_X4 FILLER_0_35_1070 ();
 FILLCELL_X2 FILLER_0_35_1079 ();
 FILLCELL_X32 FILLER_0_35_1091 ();
 FILLCELL_X16 FILLER_0_35_1123 ();
 FILLCELL_X8 FILLER_0_35_1139 ();
 FILLCELL_X1 FILLER_0_35_1147 ();
 FILLCELL_X32 FILLER_0_36_1 ();
 FILLCELL_X32 FILLER_0_36_33 ();
 FILLCELL_X32 FILLER_0_36_65 ();
 FILLCELL_X32 FILLER_0_36_97 ();
 FILLCELL_X16 FILLER_0_36_129 ();
 FILLCELL_X8 FILLER_0_36_145 ();
 FILLCELL_X4 FILLER_0_36_153 ();
 FILLCELL_X2 FILLER_0_36_157 ();
 FILLCELL_X2 FILLER_0_36_169 ();
 FILLCELL_X4 FILLER_0_36_176 ();
 FILLCELL_X1 FILLER_0_36_190 ();
 FILLCELL_X2 FILLER_0_36_216 ();
 FILLCELL_X1 FILLER_0_36_225 ();
 FILLCELL_X4 FILLER_0_36_272 ();
 FILLCELL_X1 FILLER_0_36_296 ();
 FILLCELL_X2 FILLER_0_36_385 ();
 FILLCELL_X1 FILLER_0_36_402 ();
 FILLCELL_X2 FILLER_0_36_410 ();
 FILLCELL_X1 FILLER_0_36_412 ();
 FILLCELL_X1 FILLER_0_36_423 ();
 FILLCELL_X1 FILLER_0_36_441 ();
 FILLCELL_X1 FILLER_0_36_453 ();
 FILLCELL_X1 FILLER_0_36_530 ();
 FILLCELL_X2 FILLER_0_36_629 ();
 FILLCELL_X2 FILLER_0_36_674 ();
 FILLCELL_X1 FILLER_0_36_676 ();
 FILLCELL_X2 FILLER_0_36_687 ();
 FILLCELL_X2 FILLER_0_36_702 ();
 FILLCELL_X1 FILLER_0_36_704 ();
 FILLCELL_X2 FILLER_0_36_749 ();
 FILLCELL_X2 FILLER_0_36_761 ();
 FILLCELL_X8 FILLER_0_36_780 ();
 FILLCELL_X1 FILLER_0_36_801 ();
 FILLCELL_X1 FILLER_0_36_809 ();
 FILLCELL_X2 FILLER_0_36_840 ();
 FILLCELL_X2 FILLER_0_36_893 ();
 FILLCELL_X2 FILLER_0_36_905 ();
 FILLCELL_X1 FILLER_0_36_907 ();
 FILLCELL_X2 FILLER_0_36_913 ();
 FILLCELL_X1 FILLER_0_36_915 ();
 FILLCELL_X2 FILLER_0_36_943 ();
 FILLCELL_X1 FILLER_0_36_945 ();
 FILLCELL_X2 FILLER_0_36_956 ();
 FILLCELL_X1 FILLER_0_36_982 ();
 FILLCELL_X1 FILLER_0_36_1021 ();
 FILLCELL_X1 FILLER_0_36_1037 ();
 FILLCELL_X4 FILLER_0_36_1048 ();
 FILLCELL_X2 FILLER_0_36_1052 ();
 FILLCELL_X8 FILLER_0_36_1059 ();
 FILLCELL_X32 FILLER_0_36_1083 ();
 FILLCELL_X32 FILLER_0_36_1115 ();
 FILLCELL_X1 FILLER_0_36_1147 ();
 FILLCELL_X32 FILLER_0_37_1 ();
 FILLCELL_X32 FILLER_0_37_33 ();
 FILLCELL_X32 FILLER_0_37_65 ();
 FILLCELL_X32 FILLER_0_37_97 ();
 FILLCELL_X16 FILLER_0_37_129 ();
 FILLCELL_X8 FILLER_0_37_145 ();
 FILLCELL_X4 FILLER_0_37_153 ();
 FILLCELL_X2 FILLER_0_37_157 ();
 FILLCELL_X1 FILLER_0_37_255 ();
 FILLCELL_X2 FILLER_0_37_266 ();
 FILLCELL_X1 FILLER_0_37_268 ();
 FILLCELL_X4 FILLER_0_37_279 ();
 FILLCELL_X1 FILLER_0_37_327 ();
 FILLCELL_X2 FILLER_0_37_359 ();
 FILLCELL_X2 FILLER_0_37_378 ();
 FILLCELL_X1 FILLER_0_37_380 ();
 FILLCELL_X2 FILLER_0_37_391 ();
 FILLCELL_X1 FILLER_0_37_393 ();
 FILLCELL_X1 FILLER_0_37_422 ();
 FILLCELL_X1 FILLER_0_37_450 ();
 FILLCELL_X1 FILLER_0_37_562 ();
 FILLCELL_X1 FILLER_0_37_583 ();
 FILLCELL_X2 FILLER_0_37_621 ();
 FILLCELL_X1 FILLER_0_37_662 ();
 FILLCELL_X2 FILLER_0_37_725 ();
 FILLCELL_X1 FILLER_0_37_727 ();
 FILLCELL_X1 FILLER_0_37_785 ();
 FILLCELL_X1 FILLER_0_37_790 ();
 FILLCELL_X2 FILLER_0_37_801 ();
 FILLCELL_X1 FILLER_0_37_803 ();
 FILLCELL_X4 FILLER_0_37_829 ();
 FILLCELL_X4 FILLER_0_37_843 ();
 FILLCELL_X2 FILLER_0_37_847 ();
 FILLCELL_X1 FILLER_0_37_849 ();
 FILLCELL_X1 FILLER_0_37_855 ();
 FILLCELL_X1 FILLER_0_37_866 ();
 FILLCELL_X1 FILLER_0_37_912 ();
 FILLCELL_X4 FILLER_0_37_920 ();
 FILLCELL_X2 FILLER_0_37_938 ();
 FILLCELL_X1 FILLER_0_37_940 ();
 FILLCELL_X2 FILLER_0_37_965 ();
 FILLCELL_X1 FILLER_0_37_967 ();
 FILLCELL_X4 FILLER_0_37_978 ();
 FILLCELL_X4 FILLER_0_37_999 ();
 FILLCELL_X4 FILLER_0_37_1041 ();
 FILLCELL_X2 FILLER_0_37_1065 ();
 FILLCELL_X32 FILLER_0_37_1092 ();
 FILLCELL_X16 FILLER_0_37_1124 ();
 FILLCELL_X8 FILLER_0_37_1140 ();
 FILLCELL_X32 FILLER_0_38_1 ();
 FILLCELL_X32 FILLER_0_38_33 ();
 FILLCELL_X32 FILLER_0_38_65 ();
 FILLCELL_X32 FILLER_0_38_97 ();
 FILLCELL_X16 FILLER_0_38_129 ();
 FILLCELL_X8 FILLER_0_38_145 ();
 FILLCELL_X4 FILLER_0_38_153 ();
 FILLCELL_X2 FILLER_0_38_157 ();
 FILLCELL_X1 FILLER_0_38_159 ();
 FILLCELL_X2 FILLER_0_38_170 ();
 FILLCELL_X1 FILLER_0_38_172 ();
 FILLCELL_X1 FILLER_0_38_193 ();
 FILLCELL_X1 FILLER_0_38_211 ();
 FILLCELL_X2 FILLER_0_38_243 ();
 FILLCELL_X1 FILLER_0_38_262 ();
 FILLCELL_X1 FILLER_0_38_309 ();
 FILLCELL_X1 FILLER_0_38_330 ();
 FILLCELL_X1 FILLER_0_38_358 ();
 FILLCELL_X2 FILLER_0_38_374 ();
 FILLCELL_X1 FILLER_0_38_376 ();
 FILLCELL_X2 FILLER_0_38_419 ();
 FILLCELL_X1 FILLER_0_38_431 ();
 FILLCELL_X1 FILLER_0_38_474 ();
 FILLCELL_X1 FILLER_0_38_488 ();
 FILLCELL_X2 FILLER_0_38_619 ();
 FILLCELL_X1 FILLER_0_38_729 ();
 FILLCELL_X2 FILLER_0_38_747 ();
 FILLCELL_X1 FILLER_0_38_749 ();
 FILLCELL_X2 FILLER_0_38_788 ();
 FILLCELL_X1 FILLER_0_38_790 ();
 FILLCELL_X4 FILLER_0_38_806 ();
 FILLCELL_X2 FILLER_0_38_810 ();
 FILLCELL_X1 FILLER_0_38_812 ();
 FILLCELL_X2 FILLER_0_38_816 ();
 FILLCELL_X16 FILLER_0_38_832 ();
 FILLCELL_X2 FILLER_0_38_858 ();
 FILLCELL_X4 FILLER_0_38_894 ();
 FILLCELL_X2 FILLER_0_38_898 ();
 FILLCELL_X1 FILLER_0_38_917 ();
 FILLCELL_X1 FILLER_0_38_928 ();
 FILLCELL_X1 FILLER_0_38_946 ();
 FILLCELL_X2 FILLER_0_38_964 ();
 FILLCELL_X2 FILLER_0_38_976 ();
 FILLCELL_X1 FILLER_0_38_978 ();
 FILLCELL_X2 FILLER_0_38_996 ();
 FILLCELL_X1 FILLER_0_38_998 ();
 FILLCELL_X4 FILLER_0_38_1029 ();
 FILLCELL_X2 FILLER_0_38_1033 ();
 FILLCELL_X4 FILLER_0_38_1050 ();
 FILLCELL_X1 FILLER_0_38_1054 ();
 FILLCELL_X4 FILLER_0_38_1065 ();
 FILLCELL_X4 FILLER_0_38_1074 ();
 FILLCELL_X2 FILLER_0_38_1078 ();
 FILLCELL_X1 FILLER_0_38_1080 ();
 FILLCELL_X32 FILLER_0_38_1091 ();
 FILLCELL_X16 FILLER_0_38_1123 ();
 FILLCELL_X8 FILLER_0_38_1139 ();
 FILLCELL_X1 FILLER_0_38_1147 ();
 FILLCELL_X32 FILLER_0_39_1 ();
 FILLCELL_X32 FILLER_0_39_33 ();
 FILLCELL_X32 FILLER_0_39_65 ();
 FILLCELL_X32 FILLER_0_39_97 ();
 FILLCELL_X32 FILLER_0_39_129 ();
 FILLCELL_X2 FILLER_0_39_161 ();
 FILLCELL_X1 FILLER_0_39_163 ();
 FILLCELL_X2 FILLER_0_39_179 ();
 FILLCELL_X4 FILLER_0_39_191 ();
 FILLCELL_X2 FILLER_0_39_205 ();
 FILLCELL_X1 FILLER_0_39_217 ();
 FILLCELL_X2 FILLER_0_39_235 ();
 FILLCELL_X1 FILLER_0_39_237 ();
 FILLCELL_X4 FILLER_0_39_248 ();
 FILLCELL_X2 FILLER_0_39_269 ();
 FILLCELL_X1 FILLER_0_39_271 ();
 FILLCELL_X2 FILLER_0_39_375 ();
 FILLCELL_X2 FILLER_0_39_387 ();
 FILLCELL_X1 FILLER_0_39_431 ();
 FILLCELL_X1 FILLER_0_39_465 ();
 FILLCELL_X1 FILLER_0_39_538 ();
 FILLCELL_X1 FILLER_0_39_619 ();
 FILLCELL_X2 FILLER_0_39_672 ();
 FILLCELL_X1 FILLER_0_39_711 ();
 FILLCELL_X2 FILLER_0_39_761 ();
 FILLCELL_X1 FILLER_0_39_763 ();
 FILLCELL_X8 FILLER_0_39_802 ();
 FILLCELL_X1 FILLER_0_39_816 ();
 FILLCELL_X1 FILLER_0_39_826 ();
 FILLCELL_X8 FILLER_0_39_896 ();
 FILLCELL_X1 FILLER_0_39_904 ();
 FILLCELL_X1 FILLER_0_39_936 ();
 FILLCELL_X2 FILLER_0_39_947 ();
 FILLCELL_X1 FILLER_0_39_949 ();
 FILLCELL_X2 FILLER_0_39_1030 ();
 FILLCELL_X1 FILLER_0_39_1032 ();
 FILLCELL_X1 FILLER_0_39_1052 ();
 FILLCELL_X32 FILLER_0_39_1088 ();
 FILLCELL_X16 FILLER_0_39_1120 ();
 FILLCELL_X8 FILLER_0_39_1136 ();
 FILLCELL_X4 FILLER_0_39_1144 ();
 FILLCELL_X32 FILLER_0_40_1 ();
 FILLCELL_X32 FILLER_0_40_33 ();
 FILLCELL_X32 FILLER_0_40_65 ();
 FILLCELL_X32 FILLER_0_40_97 ();
 FILLCELL_X32 FILLER_0_40_129 ();
 FILLCELL_X8 FILLER_0_40_161 ();
 FILLCELL_X2 FILLER_0_40_169 ();
 FILLCELL_X2 FILLER_0_40_200 ();
 FILLCELL_X1 FILLER_0_40_202 ();
 FILLCELL_X1 FILLER_0_40_224 ();
 FILLCELL_X2 FILLER_0_40_259 ();
 FILLCELL_X1 FILLER_0_40_261 ();
 FILLCELL_X1 FILLER_0_40_308 ();
 FILLCELL_X1 FILLER_0_40_319 ();
 FILLCELL_X1 FILLER_0_40_406 ();
 FILLCELL_X2 FILLER_0_40_417 ();
 FILLCELL_X1 FILLER_0_40_432 ();
 FILLCELL_X1 FILLER_0_40_577 ();
 FILLCELL_X1 FILLER_0_40_630 ();
 FILLCELL_X2 FILLER_0_40_654 ();
 FILLCELL_X1 FILLER_0_40_656 ();
 FILLCELL_X4 FILLER_0_40_783 ();
 FILLCELL_X2 FILLER_0_40_794 ();
 FILLCELL_X1 FILLER_0_40_796 ();
 FILLCELL_X1 FILLER_0_40_814 ();
 FILLCELL_X2 FILLER_0_40_875 ();
 FILLCELL_X2 FILLER_0_40_894 ();
 FILLCELL_X1 FILLER_0_40_900 ();
 FILLCELL_X1 FILLER_0_40_941 ();
 FILLCELL_X2 FILLER_0_40_947 ();
 FILLCELL_X2 FILLER_0_40_989 ();
 FILLCELL_X4 FILLER_0_40_1006 ();
 FILLCELL_X2 FILLER_0_40_1030 ();
 FILLCELL_X1 FILLER_0_40_1057 ();
 FILLCELL_X1 FILLER_0_40_1068 ();
 FILLCELL_X32 FILLER_0_40_1079 ();
 FILLCELL_X32 FILLER_0_40_1111 ();
 FILLCELL_X4 FILLER_0_40_1143 ();
 FILLCELL_X1 FILLER_0_40_1147 ();
 FILLCELL_X32 FILLER_0_41_1 ();
 FILLCELL_X32 FILLER_0_41_33 ();
 FILLCELL_X32 FILLER_0_41_65 ();
 FILLCELL_X32 FILLER_0_41_97 ();
 FILLCELL_X32 FILLER_0_41_129 ();
 FILLCELL_X4 FILLER_0_41_161 ();
 FILLCELL_X2 FILLER_0_41_165 ();
 FILLCELL_X1 FILLER_0_41_167 ();
 FILLCELL_X2 FILLER_0_41_212 ();
 FILLCELL_X1 FILLER_0_41_214 ();
 FILLCELL_X1 FILLER_0_41_225 ();
 FILLCELL_X1 FILLER_0_41_246 ();
 FILLCELL_X1 FILLER_0_41_254 ();
 FILLCELL_X1 FILLER_0_41_280 ();
 FILLCELL_X2 FILLER_0_41_370 ();
 FILLCELL_X2 FILLER_0_41_413 ();
 FILLCELL_X1 FILLER_0_41_422 ();
 FILLCELL_X1 FILLER_0_41_554 ();
 FILLCELL_X2 FILLER_0_41_643 ();
 FILLCELL_X1 FILLER_0_41_665 ();
 FILLCELL_X1 FILLER_0_41_679 ();
 FILLCELL_X1 FILLER_0_41_690 ();
 FILLCELL_X2 FILLER_0_41_701 ();
 FILLCELL_X1 FILLER_0_41_703 ();
 FILLCELL_X1 FILLER_0_41_780 ();
 FILLCELL_X1 FILLER_0_41_819 ();
 FILLCELL_X1 FILLER_0_41_954 ();
 FILLCELL_X2 FILLER_0_41_966 ();
 FILLCELL_X1 FILLER_0_41_968 ();
 FILLCELL_X4 FILLER_0_41_984 ();
 FILLCELL_X2 FILLER_0_41_988 ();
 FILLCELL_X1 FILLER_0_41_995 ();
 FILLCELL_X1 FILLER_0_41_1056 ();
 FILLCELL_X32 FILLER_0_41_1071 ();
 FILLCELL_X32 FILLER_0_41_1103 ();
 FILLCELL_X8 FILLER_0_41_1135 ();
 FILLCELL_X4 FILLER_0_41_1143 ();
 FILLCELL_X1 FILLER_0_41_1147 ();
 FILLCELL_X32 FILLER_0_42_1 ();
 FILLCELL_X32 FILLER_0_42_33 ();
 FILLCELL_X32 FILLER_0_42_65 ();
 FILLCELL_X32 FILLER_0_42_97 ();
 FILLCELL_X16 FILLER_0_42_129 ();
 FILLCELL_X8 FILLER_0_42_145 ();
 FILLCELL_X2 FILLER_0_42_153 ();
 FILLCELL_X1 FILLER_0_42_175 ();
 FILLCELL_X8 FILLER_0_42_186 ();
 FILLCELL_X2 FILLER_0_42_194 ();
 FILLCELL_X1 FILLER_0_42_196 ();
 FILLCELL_X1 FILLER_0_42_202 ();
 FILLCELL_X2 FILLER_0_42_213 ();
 FILLCELL_X1 FILLER_0_42_215 ();
 FILLCELL_X1 FILLER_0_42_266 ();
 FILLCELL_X4 FILLER_0_42_304 ();
 FILLCELL_X1 FILLER_0_42_318 ();
 FILLCELL_X1 FILLER_0_42_342 ();
 FILLCELL_X1 FILLER_0_42_374 ();
 FILLCELL_X4 FILLER_0_42_413 ();
 FILLCELL_X1 FILLER_0_42_542 ();
 FILLCELL_X1 FILLER_0_42_632 ();
 FILLCELL_X1 FILLER_0_42_660 ();
 FILLCELL_X1 FILLER_0_42_693 ();
 FILLCELL_X2 FILLER_0_42_714 ();
 FILLCELL_X1 FILLER_0_42_716 ();
 FILLCELL_X1 FILLER_0_42_762 ();
 FILLCELL_X2 FILLER_0_42_783 ();
 FILLCELL_X1 FILLER_0_42_785 ();
 FILLCELL_X1 FILLER_0_42_798 ();
 FILLCELL_X2 FILLER_0_42_859 ();
 FILLCELL_X2 FILLER_0_42_875 ();
 FILLCELL_X1 FILLER_0_42_894 ();
 FILLCELL_X2 FILLER_0_42_899 ();
 FILLCELL_X1 FILLER_0_42_901 ();
 FILLCELL_X16 FILLER_0_42_906 ();
 FILLCELL_X8 FILLER_0_42_922 ();
 FILLCELL_X4 FILLER_0_42_930 ();
 FILLCELL_X1 FILLER_0_42_934 ();
 FILLCELL_X2 FILLER_0_42_945 ();
 FILLCELL_X8 FILLER_0_42_957 ();
 FILLCELL_X1 FILLER_0_42_965 ();
 FILLCELL_X4 FILLER_0_42_981 ();
 FILLCELL_X2 FILLER_0_42_985 ();
 FILLCELL_X4 FILLER_0_42_1017 ();
 FILLCELL_X2 FILLER_0_42_1021 ();
 FILLCELL_X4 FILLER_0_42_1033 ();
 FILLCELL_X1 FILLER_0_42_1037 ();
 FILLCELL_X4 FILLER_0_42_1043 ();
 FILLCELL_X2 FILLER_0_42_1047 ();
 FILLCELL_X32 FILLER_0_42_1064 ();
 FILLCELL_X32 FILLER_0_42_1096 ();
 FILLCELL_X16 FILLER_0_42_1128 ();
 FILLCELL_X4 FILLER_0_42_1144 ();
 FILLCELL_X32 FILLER_0_43_1 ();
 FILLCELL_X32 FILLER_0_43_33 ();
 FILLCELL_X32 FILLER_0_43_65 ();
 FILLCELL_X32 FILLER_0_43_97 ();
 FILLCELL_X16 FILLER_0_43_129 ();
 FILLCELL_X8 FILLER_0_43_145 ();
 FILLCELL_X1 FILLER_0_43_153 ();
 FILLCELL_X1 FILLER_0_43_169 ();
 FILLCELL_X1 FILLER_0_43_180 ();
 FILLCELL_X4 FILLER_0_43_195 ();
 FILLCELL_X1 FILLER_0_43_199 ();
 FILLCELL_X2 FILLER_0_43_217 ();
 FILLCELL_X1 FILLER_0_43_270 ();
 FILLCELL_X4 FILLER_0_43_304 ();
 FILLCELL_X1 FILLER_0_43_325 ();
 FILLCELL_X1 FILLER_0_43_404 ();
 FILLCELL_X1 FILLER_0_43_543 ();
 FILLCELL_X2 FILLER_0_43_638 ();
 FILLCELL_X2 FILLER_0_43_650 ();
 FILLCELL_X1 FILLER_0_43_652 ();
 FILLCELL_X1 FILLER_0_43_690 ();
 FILLCELL_X2 FILLER_0_43_708 ();
 FILLCELL_X1 FILLER_0_43_710 ();
 FILLCELL_X1 FILLER_0_43_814 ();
 FILLCELL_X1 FILLER_0_43_819 ();
 FILLCELL_X1 FILLER_0_43_861 ();
 FILLCELL_X1 FILLER_0_43_890 ();
 FILLCELL_X2 FILLER_0_43_908 ();
 FILLCELL_X8 FILLER_0_43_917 ();
 FILLCELL_X2 FILLER_0_43_925 ();
 FILLCELL_X1 FILLER_0_43_927 ();
 FILLCELL_X8 FILLER_0_43_933 ();
 FILLCELL_X4 FILLER_0_43_941 ();
 FILLCELL_X2 FILLER_0_43_945 ();
 FILLCELL_X4 FILLER_0_43_954 ();
 FILLCELL_X1 FILLER_0_43_958 ();
 FILLCELL_X8 FILLER_0_43_974 ();
 FILLCELL_X2 FILLER_0_43_982 ();
 FILLCELL_X8 FILLER_0_43_991 ();
 FILLCELL_X2 FILLER_0_43_999 ();
 FILLCELL_X1 FILLER_0_43_1001 ();
 FILLCELL_X2 FILLER_0_43_1007 ();
 FILLCELL_X1 FILLER_0_43_1009 ();
 FILLCELL_X32 FILLER_0_43_1015 ();
 FILLCELL_X32 FILLER_0_43_1047 ();
 FILLCELL_X32 FILLER_0_43_1079 ();
 FILLCELL_X32 FILLER_0_43_1111 ();
 FILLCELL_X4 FILLER_0_43_1143 ();
 FILLCELL_X1 FILLER_0_43_1147 ();
 FILLCELL_X32 FILLER_0_44_1 ();
 FILLCELL_X32 FILLER_0_44_33 ();
 FILLCELL_X32 FILLER_0_44_65 ();
 FILLCELL_X32 FILLER_0_44_97 ();
 FILLCELL_X32 FILLER_0_44_129 ();
 FILLCELL_X4 FILLER_0_44_161 ();
 FILLCELL_X1 FILLER_0_44_165 ();
 FILLCELL_X4 FILLER_0_44_176 ();
 FILLCELL_X2 FILLER_0_44_189 ();
 FILLCELL_X8 FILLER_0_44_201 ();
 FILLCELL_X1 FILLER_0_44_209 ();
 FILLCELL_X8 FILLER_0_44_215 ();
 FILLCELL_X1 FILLER_0_44_223 ();
 FILLCELL_X1 FILLER_0_44_234 ();
 FILLCELL_X1 FILLER_0_44_240 ();
 FILLCELL_X1 FILLER_0_44_309 ();
 FILLCELL_X4 FILLER_0_44_403 ();
 FILLCELL_X2 FILLER_0_44_407 ();
 FILLCELL_X1 FILLER_0_44_543 ();
 FILLCELL_X1 FILLER_0_44_586 ();
 FILLCELL_X1 FILLER_0_44_607 ();
 FILLCELL_X1 FILLER_0_44_630 ();
 FILLCELL_X2 FILLER_0_44_632 ();
 FILLCELL_X1 FILLER_0_44_634 ();
 FILLCELL_X1 FILLER_0_44_856 ();
 FILLCELL_X1 FILLER_0_44_865 ();
 FILLCELL_X2 FILLER_0_44_872 ();
 FILLCELL_X1 FILLER_0_44_899 ();
 FILLCELL_X1 FILLER_0_44_910 ();
 FILLCELL_X2 FILLER_0_44_965 ();
 FILLCELL_X4 FILLER_0_44_1022 ();
 FILLCELL_X2 FILLER_0_44_1026 ();
 FILLCELL_X1 FILLER_0_44_1028 ();
 FILLCELL_X8 FILLER_0_44_1034 ();
 FILLCELL_X1 FILLER_0_44_1042 ();
 FILLCELL_X32 FILLER_0_44_1073 ();
 FILLCELL_X32 FILLER_0_44_1105 ();
 FILLCELL_X8 FILLER_0_44_1137 ();
 FILLCELL_X2 FILLER_0_44_1145 ();
 FILLCELL_X1 FILLER_0_44_1147 ();
 FILLCELL_X32 FILLER_0_45_1 ();
 FILLCELL_X32 FILLER_0_45_33 ();
 FILLCELL_X32 FILLER_0_45_65 ();
 FILLCELL_X32 FILLER_0_45_97 ();
 FILLCELL_X16 FILLER_0_45_129 ();
 FILLCELL_X8 FILLER_0_45_145 ();
 FILLCELL_X1 FILLER_0_45_153 ();
 FILLCELL_X2 FILLER_0_45_179 ();
 FILLCELL_X1 FILLER_0_45_181 ();
 FILLCELL_X16 FILLER_0_45_192 ();
 FILLCELL_X4 FILLER_0_45_208 ();
 FILLCELL_X1 FILLER_0_45_212 ();
 FILLCELL_X4 FILLER_0_45_223 ();
 FILLCELL_X2 FILLER_0_45_227 ();
 FILLCELL_X1 FILLER_0_45_233 ();
 FILLCELL_X2 FILLER_0_45_239 ();
 FILLCELL_X2 FILLER_0_45_279 ();
 FILLCELL_X2 FILLER_0_45_290 ();
 FILLCELL_X2 FILLER_0_45_302 ();
 FILLCELL_X4 FILLER_0_45_316 ();
 FILLCELL_X2 FILLER_0_45_344 ();
 FILLCELL_X1 FILLER_0_45_452 ();
 FILLCELL_X2 FILLER_0_45_460 ();
 FILLCELL_X1 FILLER_0_45_562 ();
 FILLCELL_X2 FILLER_0_45_611 ();
 FILLCELL_X2 FILLER_0_45_681 ();
 FILLCELL_X1 FILLER_0_45_683 ();
 FILLCELL_X1 FILLER_0_45_694 ();
 FILLCELL_X2 FILLER_0_45_712 ();
 FILLCELL_X1 FILLER_0_45_807 ();
 FILLCELL_X2 FILLER_0_45_838 ();
 FILLCELL_X2 FILLER_0_45_880 ();
 FILLCELL_X1 FILLER_0_45_889 ();
 FILLCELL_X4 FILLER_0_45_915 ();
 FILLCELL_X2 FILLER_0_45_929 ();
 FILLCELL_X1 FILLER_0_45_931 ();
 FILLCELL_X2 FILLER_0_45_947 ();
 FILLCELL_X1 FILLER_0_45_949 ();
 FILLCELL_X2 FILLER_0_45_960 ();
 FILLCELL_X1 FILLER_0_45_962 ();
 FILLCELL_X2 FILLER_0_45_1015 ();
 FILLCELL_X32 FILLER_0_45_1077 ();
 FILLCELL_X32 FILLER_0_45_1109 ();
 FILLCELL_X4 FILLER_0_45_1141 ();
 FILLCELL_X2 FILLER_0_45_1145 ();
 FILLCELL_X1 FILLER_0_45_1147 ();
 FILLCELL_X32 FILLER_0_46_1 ();
 FILLCELL_X32 FILLER_0_46_33 ();
 FILLCELL_X32 FILLER_0_46_65 ();
 FILLCELL_X32 FILLER_0_46_97 ();
 FILLCELL_X32 FILLER_0_46_129 ();
 FILLCELL_X4 FILLER_0_46_161 ();
 FILLCELL_X2 FILLER_0_46_165 ();
 FILLCELL_X2 FILLER_0_46_177 ();
 FILLCELL_X1 FILLER_0_46_179 ();
 FILLCELL_X1 FILLER_0_46_209 ();
 FILLCELL_X4 FILLER_0_46_235 ();
 FILLCELL_X1 FILLER_0_46_249 ();
 FILLCELL_X1 FILLER_0_46_259 ();
 FILLCELL_X1 FILLER_0_46_294 ();
 FILLCELL_X1 FILLER_0_46_305 ();
 FILLCELL_X1 FILLER_0_46_356 ();
 FILLCELL_X1 FILLER_0_46_447 ();
 FILLCELL_X2 FILLER_0_46_628 ();
 FILLCELL_X1 FILLER_0_46_630 ();
 FILLCELL_X4 FILLER_0_46_662 ();
 FILLCELL_X2 FILLER_0_46_693 ();
 FILLCELL_X1 FILLER_0_46_724 ();
 FILLCELL_X1 FILLER_0_46_754 ();
 FILLCELL_X2 FILLER_0_46_802 ();
 FILLCELL_X1 FILLER_0_46_846 ();
 FILLCELL_X2 FILLER_0_46_920 ();
 FILLCELL_X1 FILLER_0_46_922 ();
 FILLCELL_X2 FILLER_0_46_979 ();
 FILLCELL_X4 FILLER_0_46_1016 ();
 FILLCELL_X1 FILLER_0_46_1035 ();
 FILLCELL_X32 FILLER_0_46_1080 ();
 FILLCELL_X32 FILLER_0_46_1112 ();
 FILLCELL_X4 FILLER_0_46_1144 ();
 FILLCELL_X32 FILLER_0_47_1 ();
 FILLCELL_X32 FILLER_0_47_33 ();
 FILLCELL_X32 FILLER_0_47_65 ();
 FILLCELL_X32 FILLER_0_47_97 ();
 FILLCELL_X32 FILLER_0_47_129 ();
 FILLCELL_X4 FILLER_0_47_161 ();
 FILLCELL_X1 FILLER_0_47_165 ();
 FILLCELL_X1 FILLER_0_47_176 ();
 FILLCELL_X2 FILLER_0_47_187 ();
 FILLCELL_X1 FILLER_0_47_189 ();
 FILLCELL_X1 FILLER_0_47_200 ();
 FILLCELL_X4 FILLER_0_47_206 ();
 FILLCELL_X2 FILLER_0_47_210 ();
 FILLCELL_X1 FILLER_0_47_212 ();
 FILLCELL_X2 FILLER_0_47_217 ();
 FILLCELL_X8 FILLER_0_47_243 ();
 FILLCELL_X2 FILLER_0_47_251 ();
 FILLCELL_X1 FILLER_0_47_253 ();
 FILLCELL_X2 FILLER_0_47_264 ();
 FILLCELL_X4 FILLER_0_47_293 ();
 FILLCELL_X1 FILLER_0_47_334 ();
 FILLCELL_X1 FILLER_0_47_348 ();
 FILLCELL_X1 FILLER_0_47_358 ();
 FILLCELL_X1 FILLER_0_47_569 ();
 FILLCELL_X4 FILLER_0_47_638 ();
 FILLCELL_X4 FILLER_0_47_659 ();
 FILLCELL_X1 FILLER_0_47_678 ();
 FILLCELL_X2 FILLER_0_47_703 ();
 FILLCELL_X2 FILLER_0_47_720 ();
 FILLCELL_X1 FILLER_0_47_786 ();
 FILLCELL_X2 FILLER_0_47_799 ();
 FILLCELL_X1 FILLER_0_47_828 ();
 FILLCELL_X2 FILLER_0_47_897 ();
 FILLCELL_X1 FILLER_0_47_899 ();
 FILLCELL_X1 FILLER_0_47_925 ();
 FILLCELL_X1 FILLER_0_47_959 ();
 FILLCELL_X1 FILLER_0_47_977 ();
 FILLCELL_X4 FILLER_0_47_1062 ();
 FILLCELL_X1 FILLER_0_47_1066 ();
 FILLCELL_X32 FILLER_0_47_1077 ();
 FILLCELL_X32 FILLER_0_47_1109 ();
 FILLCELL_X4 FILLER_0_47_1141 ();
 FILLCELL_X2 FILLER_0_47_1145 ();
 FILLCELL_X1 FILLER_0_47_1147 ();
 FILLCELL_X32 FILLER_0_48_1 ();
 FILLCELL_X32 FILLER_0_48_33 ();
 FILLCELL_X32 FILLER_0_48_65 ();
 FILLCELL_X32 FILLER_0_48_97 ();
 FILLCELL_X16 FILLER_0_48_129 ();
 FILLCELL_X8 FILLER_0_48_145 ();
 FILLCELL_X4 FILLER_0_48_153 ();
 FILLCELL_X2 FILLER_0_48_157 ();
 FILLCELL_X4 FILLER_0_48_193 ();
 FILLCELL_X16 FILLER_0_48_227 ();
 FILLCELL_X8 FILLER_0_48_243 ();
 FILLCELL_X2 FILLER_0_48_281 ();
 FILLCELL_X1 FILLER_0_48_283 ();
 FILLCELL_X1 FILLER_0_48_313 ();
 FILLCELL_X1 FILLER_0_48_349 ();
 FILLCELL_X1 FILLER_0_48_370 ();
 FILLCELL_X1 FILLER_0_48_385 ();
 FILLCELL_X1 FILLER_0_48_530 ();
 FILLCELL_X1 FILLER_0_48_620 ();
 FILLCELL_X2 FILLER_0_48_659 ();
 FILLCELL_X1 FILLER_0_48_661 ();
 FILLCELL_X2 FILLER_0_48_697 ();
 FILLCELL_X1 FILLER_0_48_699 ();
 FILLCELL_X2 FILLER_0_48_723 ();
 FILLCELL_X1 FILLER_0_48_725 ();
 FILLCELL_X2 FILLER_0_48_758 ();
 FILLCELL_X1 FILLER_0_48_867 ();
 FILLCELL_X2 FILLER_0_48_897 ();
 FILLCELL_X1 FILLER_0_48_909 ();
 FILLCELL_X4 FILLER_0_48_931 ();
 FILLCELL_X1 FILLER_0_48_952 ();
 FILLCELL_X1 FILLER_0_48_963 ();
 FILLCELL_X4 FILLER_0_48_1019 ();
 FILLCELL_X1 FILLER_0_48_1033 ();
 FILLCELL_X1 FILLER_0_48_1054 ();
 FILLCELL_X32 FILLER_0_48_1070 ();
 FILLCELL_X32 FILLER_0_48_1102 ();
 FILLCELL_X8 FILLER_0_48_1134 ();
 FILLCELL_X4 FILLER_0_48_1142 ();
 FILLCELL_X2 FILLER_0_48_1146 ();
 FILLCELL_X32 FILLER_0_49_1 ();
 FILLCELL_X32 FILLER_0_49_33 ();
 FILLCELL_X32 FILLER_0_49_65 ();
 FILLCELL_X32 FILLER_0_49_97 ();
 FILLCELL_X32 FILLER_0_49_129 ();
 FILLCELL_X32 FILLER_0_49_161 ();
 FILLCELL_X2 FILLER_0_49_193 ();
 FILLCELL_X32 FILLER_0_49_205 ();
 FILLCELL_X2 FILLER_0_49_237 ();
 FILLCELL_X1 FILLER_0_49_239 ();
 FILLCELL_X4 FILLER_0_49_301 ();
 FILLCELL_X1 FILLER_0_49_310 ();
 FILLCELL_X1 FILLER_0_49_334 ();
 FILLCELL_X1 FILLER_0_49_395 ();
 FILLCELL_X1 FILLER_0_49_428 ();
 FILLCELL_X2 FILLER_0_49_484 ();
 FILLCELL_X1 FILLER_0_49_606 ();
 FILLCELL_X2 FILLER_0_49_636 ();
 FILLCELL_X1 FILLER_0_49_638 ();
 FILLCELL_X1 FILLER_0_49_671 ();
 FILLCELL_X1 FILLER_0_49_687 ();
 FILLCELL_X2 FILLER_0_49_718 ();
 FILLCELL_X1 FILLER_0_49_720 ();
 FILLCELL_X2 FILLER_0_49_832 ();
 FILLCELL_X2 FILLER_0_49_858 ();
 FILLCELL_X1 FILLER_0_49_870 ();
 FILLCELL_X2 FILLER_0_49_886 ();
 FILLCELL_X4 FILLER_0_49_903 ();
 FILLCELL_X1 FILLER_0_49_914 ();
 FILLCELL_X1 FILLER_0_49_930 ();
 FILLCELL_X2 FILLER_0_49_963 ();
 FILLCELL_X4 FILLER_0_49_1034 ();
 FILLCELL_X1 FILLER_0_49_1048 ();
 FILLCELL_X4 FILLER_0_49_1074 ();
 FILLCELL_X2 FILLER_0_49_1078 ();
 FILLCELL_X8 FILLER_0_49_1090 ();
 FILLCELL_X4 FILLER_0_49_1098 ();
 FILLCELL_X2 FILLER_0_49_1102 ();
 FILLCELL_X1 FILLER_0_49_1104 ();
 FILLCELL_X16 FILLER_0_49_1112 ();
 FILLCELL_X8 FILLER_0_49_1135 ();
 FILLCELL_X4 FILLER_0_49_1143 ();
 FILLCELL_X1 FILLER_0_49_1147 ();
 FILLCELL_X32 FILLER_0_50_1 ();
 FILLCELL_X32 FILLER_0_50_33 ();
 FILLCELL_X32 FILLER_0_50_65 ();
 FILLCELL_X32 FILLER_0_50_97 ();
 FILLCELL_X32 FILLER_0_50_129 ();
 FILLCELL_X16 FILLER_0_50_161 ();
 FILLCELL_X4 FILLER_0_50_177 ();
 FILLCELL_X1 FILLER_0_50_181 ();
 FILLCELL_X4 FILLER_0_50_187 ();
 FILLCELL_X4 FILLER_0_50_206 ();
 FILLCELL_X4 FILLER_0_50_222 ();
 FILLCELL_X1 FILLER_0_50_287 ();
 FILLCELL_X1 FILLER_0_50_298 ();
 FILLCELL_X1 FILLER_0_50_320 ();
 FILLCELL_X2 FILLER_0_50_345 ();
 FILLCELL_X1 FILLER_0_50_385 ();
 FILLCELL_X2 FILLER_0_50_483 ();
 FILLCELL_X2 FILLER_0_50_628 ();
 FILLCELL_X1 FILLER_0_50_630 ();
 FILLCELL_X2 FILLER_0_50_644 ();
 FILLCELL_X1 FILLER_0_50_646 ();
 FILLCELL_X4 FILLER_0_50_667 ();
 FILLCELL_X1 FILLER_0_50_682 ();
 FILLCELL_X1 FILLER_0_50_697 ();
 FILLCELL_X2 FILLER_0_50_708 ();
 FILLCELL_X1 FILLER_0_50_813 ();
 FILLCELL_X1 FILLER_0_50_825 ();
 FILLCELL_X4 FILLER_0_50_882 ();
 FILLCELL_X2 FILLER_0_50_930 ();
 FILLCELL_X1 FILLER_0_50_932 ();
 FILLCELL_X2 FILLER_0_50_954 ();
 FILLCELL_X1 FILLER_0_50_956 ();
 FILLCELL_X2 FILLER_0_50_981 ();
 FILLCELL_X1 FILLER_0_50_1002 ();
 FILLCELL_X2 FILLER_0_50_1043 ();
 FILLCELL_X2 FILLER_0_50_1050 ();
 FILLCELL_X32 FILLER_0_50_1072 ();
 FILLCELL_X2 FILLER_0_50_1104 ();
 FILLCELL_X1 FILLER_0_50_1106 ();
 FILLCELL_X32 FILLER_0_50_1114 ();
 FILLCELL_X2 FILLER_0_50_1146 ();
 FILLCELL_X32 FILLER_0_51_1 ();
 FILLCELL_X32 FILLER_0_51_33 ();
 FILLCELL_X32 FILLER_0_51_65 ();
 FILLCELL_X32 FILLER_0_51_97 ();
 FILLCELL_X32 FILLER_0_51_129 ();
 FILLCELL_X2 FILLER_0_51_161 ();
 FILLCELL_X1 FILLER_0_51_202 ();
 FILLCELL_X4 FILLER_0_51_232 ();
 FILLCELL_X2 FILLER_0_51_253 ();
 FILLCELL_X1 FILLER_0_51_255 ();
 FILLCELL_X2 FILLER_0_51_266 ();
 FILLCELL_X1 FILLER_0_51_285 ();
 FILLCELL_X2 FILLER_0_51_296 ();
 FILLCELL_X1 FILLER_0_51_298 ();
 FILLCELL_X2 FILLER_0_51_309 ();
 FILLCELL_X1 FILLER_0_51_311 ();
 FILLCELL_X1 FILLER_0_51_361 ();
 FILLCELL_X8 FILLER_0_51_369 ();
 FILLCELL_X2 FILLER_0_51_387 ();
 FILLCELL_X2 FILLER_0_51_429 ();
 FILLCELL_X2 FILLER_0_51_457 ();
 FILLCELL_X1 FILLER_0_51_459 ();
 FILLCELL_X1 FILLER_0_51_555 ();
 FILLCELL_X1 FILLER_0_51_629 ();
 FILLCELL_X2 FILLER_0_51_652 ();
 FILLCELL_X1 FILLER_0_51_654 ();
 FILLCELL_X2 FILLER_0_51_680 ();
 FILLCELL_X1 FILLER_0_51_682 ();
 FILLCELL_X2 FILLER_0_51_876 ();
 FILLCELL_X1 FILLER_0_51_878 ();
 FILLCELL_X2 FILLER_0_51_884 ();
 FILLCELL_X1 FILLER_0_51_896 ();
 FILLCELL_X2 FILLER_0_51_907 ();
 FILLCELL_X1 FILLER_0_51_909 ();
 FILLCELL_X2 FILLER_0_51_917 ();
 FILLCELL_X2 FILLER_0_51_929 ();
 FILLCELL_X1 FILLER_0_51_975 ();
 FILLCELL_X4 FILLER_0_51_1003 ();
 FILLCELL_X2 FILLER_0_51_1062 ();
 FILLCELL_X32 FILLER_0_51_1074 ();
 FILLCELL_X8 FILLER_0_51_1106 ();
 FILLCELL_X16 FILLER_0_51_1128 ();
 FILLCELL_X4 FILLER_0_51_1144 ();
 FILLCELL_X32 FILLER_0_52_1 ();
 FILLCELL_X32 FILLER_0_52_33 ();
 FILLCELL_X32 FILLER_0_52_65 ();
 FILLCELL_X32 FILLER_0_52_97 ();
 FILLCELL_X32 FILLER_0_52_129 ();
 FILLCELL_X2 FILLER_0_52_161 ();
 FILLCELL_X2 FILLER_0_52_173 ();
 FILLCELL_X1 FILLER_0_52_175 ();
 FILLCELL_X2 FILLER_0_52_181 ();
 FILLCELL_X4 FILLER_0_52_193 ();
 FILLCELL_X1 FILLER_0_52_214 ();
 FILLCELL_X4 FILLER_0_52_271 ();
 FILLCELL_X4 FILLER_0_52_282 ();
 FILLCELL_X4 FILLER_0_52_378 ();
 FILLCELL_X2 FILLER_0_52_382 ();
 FILLCELL_X2 FILLER_0_52_405 ();
 FILLCELL_X1 FILLER_0_52_407 ();
 FILLCELL_X1 FILLER_0_52_413 ();
 FILLCELL_X2 FILLER_0_52_424 ();
 FILLCELL_X1 FILLER_0_52_495 ();
 FILLCELL_X1 FILLER_0_52_615 ();
 FILLCELL_X1 FILLER_0_52_632 ();
 FILLCELL_X2 FILLER_0_52_643 ();
 FILLCELL_X4 FILLER_0_52_655 ();
 FILLCELL_X2 FILLER_0_52_674 ();
 FILLCELL_X2 FILLER_0_52_686 ();
 FILLCELL_X1 FILLER_0_52_688 ();
 FILLCELL_X2 FILLER_0_52_708 ();
 FILLCELL_X1 FILLER_0_52_730 ();
 FILLCELL_X2 FILLER_0_52_764 ();
 FILLCELL_X1 FILLER_0_52_790 ();
 FILLCELL_X1 FILLER_0_52_843 ();
 FILLCELL_X2 FILLER_0_52_881 ();
 FILLCELL_X1 FILLER_0_52_883 ();
 FILLCELL_X4 FILLER_0_52_960 ();
 FILLCELL_X2 FILLER_0_52_974 ();
 FILLCELL_X2 FILLER_0_52_1000 ();
 FILLCELL_X1 FILLER_0_52_1002 ();
 FILLCELL_X2 FILLER_0_52_1027 ();
 FILLCELL_X1 FILLER_0_52_1029 ();
 FILLCELL_X2 FILLER_0_52_1050 ();
 FILLCELL_X1 FILLER_0_52_1052 ();
 FILLCELL_X4 FILLER_0_52_1063 ();
 FILLCELL_X32 FILLER_0_52_1077 ();
 FILLCELL_X32 FILLER_0_52_1109 ();
 FILLCELL_X4 FILLER_0_52_1141 ();
 FILLCELL_X2 FILLER_0_52_1145 ();
 FILLCELL_X1 FILLER_0_52_1147 ();
 FILLCELL_X32 FILLER_0_53_1 ();
 FILLCELL_X32 FILLER_0_53_33 ();
 FILLCELL_X32 FILLER_0_53_65 ();
 FILLCELL_X32 FILLER_0_53_97 ();
 FILLCELL_X32 FILLER_0_53_129 ();
 FILLCELL_X4 FILLER_0_53_161 ();
 FILLCELL_X1 FILLER_0_53_165 ();
 FILLCELL_X1 FILLER_0_53_196 ();
 FILLCELL_X2 FILLER_0_53_212 ();
 FILLCELL_X2 FILLER_0_53_261 ();
 FILLCELL_X1 FILLER_0_53_263 ();
 FILLCELL_X2 FILLER_0_53_281 ();
 FILLCELL_X1 FILLER_0_53_382 ();
 FILLCELL_X1 FILLER_0_53_387 ();
 FILLCELL_X1 FILLER_0_53_398 ();
 FILLCELL_X1 FILLER_0_53_458 ();
 FILLCELL_X2 FILLER_0_53_474 ();
 FILLCELL_X1 FILLER_0_53_546 ();
 FILLCELL_X1 FILLER_0_53_583 ();
 FILLCELL_X4 FILLER_0_53_600 ();
 FILLCELL_X2 FILLER_0_53_614 ();
 FILLCELL_X1 FILLER_0_53_685 ();
 FILLCELL_X8 FILLER_0_53_742 ();
 FILLCELL_X4 FILLER_0_53_750 ();
 FILLCELL_X2 FILLER_0_53_754 ();
 FILLCELL_X2 FILLER_0_53_798 ();
 FILLCELL_X2 FILLER_0_53_851 ();
 FILLCELL_X1 FILLER_0_53_853 ();
 FILLCELL_X1 FILLER_0_53_864 ();
 FILLCELL_X2 FILLER_0_53_889 ();
 FILLCELL_X2 FILLER_0_53_923 ();
 FILLCELL_X1 FILLER_0_53_925 ();
 FILLCELL_X4 FILLER_0_53_993 ();
 FILLCELL_X1 FILLER_0_53_1032 ();
 FILLCELL_X4 FILLER_0_53_1048 ();
 FILLCELL_X4 FILLER_0_53_1062 ();
 FILLCELL_X2 FILLER_0_53_1075 ();
 FILLCELL_X1 FILLER_0_53_1077 ();
 FILLCELL_X32 FILLER_0_53_1088 ();
 FILLCELL_X16 FILLER_0_53_1120 ();
 FILLCELL_X8 FILLER_0_53_1136 ();
 FILLCELL_X4 FILLER_0_53_1144 ();
 FILLCELL_X32 FILLER_0_54_1 ();
 FILLCELL_X32 FILLER_0_54_33 ();
 FILLCELL_X32 FILLER_0_54_65 ();
 FILLCELL_X32 FILLER_0_54_97 ();
 FILLCELL_X32 FILLER_0_54_129 ();
 FILLCELL_X8 FILLER_0_54_161 ();
 FILLCELL_X4 FILLER_0_54_261 ();
 FILLCELL_X4 FILLER_0_54_308 ();
 FILLCELL_X1 FILLER_0_54_336 ();
 FILLCELL_X4 FILLER_0_54_393 ();
 FILLCELL_X8 FILLER_0_54_407 ();
 FILLCELL_X2 FILLER_0_54_415 ();
 FILLCELL_X1 FILLER_0_54_417 ();
 FILLCELL_X2 FILLER_0_54_443 ();
 FILLCELL_X1 FILLER_0_54_445 ();
 FILLCELL_X1 FILLER_0_54_537 ();
 FILLCELL_X1 FILLER_0_54_593 ();
 FILLCELL_X1 FILLER_0_54_632 ();
 FILLCELL_X1 FILLER_0_54_643 ();
 FILLCELL_X1 FILLER_0_54_649 ();
 FILLCELL_X2 FILLER_0_54_660 ();
 FILLCELL_X2 FILLER_0_54_667 ();
 FILLCELL_X1 FILLER_0_54_669 ();
 FILLCELL_X1 FILLER_0_54_705 ();
 FILLCELL_X4 FILLER_0_54_713 ();
 FILLCELL_X2 FILLER_0_54_717 ();
 FILLCELL_X1 FILLER_0_54_719 ();
 FILLCELL_X4 FILLER_0_54_725 ();
 FILLCELL_X1 FILLER_0_54_729 ();
 FILLCELL_X2 FILLER_0_54_744 ();
 FILLCELL_X2 FILLER_0_54_756 ();
 FILLCELL_X2 FILLER_0_54_768 ();
 FILLCELL_X1 FILLER_0_54_770 ();
 FILLCELL_X1 FILLER_0_54_817 ();
 FILLCELL_X2 FILLER_0_54_841 ();
 FILLCELL_X4 FILLER_0_54_885 ();
 FILLCELL_X2 FILLER_0_54_928 ();
 FILLCELL_X4 FILLER_0_54_961 ();
 FILLCELL_X2 FILLER_0_54_1049 ();
 FILLCELL_X1 FILLER_0_54_1066 ();
 FILLCELL_X1 FILLER_0_54_1077 ();
 FILLCELL_X32 FILLER_0_54_1088 ();
 FILLCELL_X16 FILLER_0_54_1120 ();
 FILLCELL_X8 FILLER_0_54_1136 ();
 FILLCELL_X4 FILLER_0_54_1144 ();
 FILLCELL_X32 FILLER_0_55_1 ();
 FILLCELL_X32 FILLER_0_55_33 ();
 FILLCELL_X32 FILLER_0_55_65 ();
 FILLCELL_X32 FILLER_0_55_97 ();
 FILLCELL_X32 FILLER_0_55_129 ();
 FILLCELL_X2 FILLER_0_55_161 ();
 FILLCELL_X1 FILLER_0_55_163 ();
 FILLCELL_X2 FILLER_0_55_197 ();
 FILLCELL_X2 FILLER_0_55_223 ();
 FILLCELL_X1 FILLER_0_55_281 ();
 FILLCELL_X2 FILLER_0_55_379 ();
 FILLCELL_X1 FILLER_0_55_381 ();
 FILLCELL_X2 FILLER_0_55_391 ();
 FILLCELL_X4 FILLER_0_55_403 ();
 FILLCELL_X1 FILLER_0_55_407 ();
 FILLCELL_X4 FILLER_0_55_410 ();
 FILLCELL_X2 FILLER_0_55_414 ();
 FILLCELL_X1 FILLER_0_55_416 ();
 FILLCELL_X2 FILLER_0_55_429 ();
 FILLCELL_X1 FILLER_0_55_441 ();
 FILLCELL_X2 FILLER_0_55_466 ();
 FILLCELL_X1 FILLER_0_55_468 ();
 FILLCELL_X4 FILLER_0_55_486 ();
 FILLCELL_X1 FILLER_0_55_540 ();
 FILLCELL_X1 FILLER_0_55_589 ();
 FILLCELL_X2 FILLER_0_55_601 ();
 FILLCELL_X1 FILLER_0_55_603 ();
 FILLCELL_X1 FILLER_0_55_634 ();
 FILLCELL_X4 FILLER_0_55_653 ();
 FILLCELL_X2 FILLER_0_55_657 ();
 FILLCELL_X1 FILLER_0_55_664 ();
 FILLCELL_X2 FILLER_0_55_675 ();
 FILLCELL_X2 FILLER_0_55_696 ();
 FILLCELL_X1 FILLER_0_55_698 ();
 FILLCELL_X8 FILLER_0_55_706 ();
 FILLCELL_X4 FILLER_0_55_732 ();
 FILLCELL_X1 FILLER_0_55_746 ();
 FILLCELL_X8 FILLER_0_55_751 ();
 FILLCELL_X2 FILLER_0_55_759 ();
 FILLCELL_X2 FILLER_0_55_765 ();
 FILLCELL_X2 FILLER_0_55_781 ();
 FILLCELL_X1 FILLER_0_55_843 ();
 FILLCELL_X1 FILLER_0_55_917 ();
 FILLCELL_X1 FILLER_0_55_933 ();
 FILLCELL_X2 FILLER_0_55_944 ();
 FILLCELL_X1 FILLER_0_55_946 ();
 FILLCELL_X2 FILLER_0_55_969 ();
 FILLCELL_X2 FILLER_0_55_998 ();
 FILLCELL_X1 FILLER_0_55_1000 ();
 FILLCELL_X2 FILLER_0_55_1056 ();
 FILLCELL_X1 FILLER_0_55_1058 ();
 FILLCELL_X32 FILLER_0_55_1088 ();
 FILLCELL_X16 FILLER_0_55_1120 ();
 FILLCELL_X8 FILLER_0_55_1136 ();
 FILLCELL_X4 FILLER_0_55_1144 ();
 FILLCELL_X32 FILLER_0_56_1 ();
 FILLCELL_X32 FILLER_0_56_33 ();
 FILLCELL_X32 FILLER_0_56_65 ();
 FILLCELL_X32 FILLER_0_56_97 ();
 FILLCELL_X32 FILLER_0_56_129 ();
 FILLCELL_X1 FILLER_0_56_201 ();
 FILLCELL_X1 FILLER_0_56_229 ();
 FILLCELL_X2 FILLER_0_56_258 ();
 FILLCELL_X1 FILLER_0_56_260 ();
 FILLCELL_X2 FILLER_0_56_271 ();
 FILLCELL_X1 FILLER_0_56_273 ();
 FILLCELL_X2 FILLER_0_56_298 ();
 FILLCELL_X1 FILLER_0_56_300 ();
 FILLCELL_X2 FILLER_0_56_381 ();
 FILLCELL_X2 FILLER_0_56_387 ();
 FILLCELL_X1 FILLER_0_56_389 ();
 FILLCELL_X1 FILLER_0_56_438 ();
 FILLCELL_X2 FILLER_0_56_452 ();
 FILLCELL_X2 FILLER_0_56_460 ();
 FILLCELL_X1 FILLER_0_56_462 ();
 FILLCELL_X1 FILLER_0_56_486 ();
 FILLCELL_X2 FILLER_0_56_497 ();
 FILLCELL_X1 FILLER_0_56_595 ();
 FILLCELL_X2 FILLER_0_56_640 ();
 FILLCELL_X16 FILLER_0_56_684 ();
 FILLCELL_X2 FILLER_0_56_714 ();
 FILLCELL_X1 FILLER_0_56_716 ();
 FILLCELL_X1 FILLER_0_56_750 ();
 FILLCELL_X1 FILLER_0_56_766 ();
 FILLCELL_X2 FILLER_0_56_771 ();
 FILLCELL_X1 FILLER_0_56_799 ();
 FILLCELL_X1 FILLER_0_56_807 ();
 FILLCELL_X1 FILLER_0_56_832 ();
 FILLCELL_X1 FILLER_0_56_843 ();
 FILLCELL_X2 FILLER_0_56_870 ();
 FILLCELL_X2 FILLER_0_56_877 ();
 FILLCELL_X1 FILLER_0_56_879 ();
 FILLCELL_X1 FILLER_0_56_890 ();
 FILLCELL_X2 FILLER_0_56_904 ();
 FILLCELL_X1 FILLER_0_56_906 ();
 FILLCELL_X2 FILLER_0_56_980 ();
 FILLCELL_X1 FILLER_0_56_982 ();
 FILLCELL_X2 FILLER_0_56_1032 ();
 FILLCELL_X1 FILLER_0_56_1034 ();
 FILLCELL_X1 FILLER_0_56_1045 ();
 FILLCELL_X32 FILLER_0_56_1076 ();
 FILLCELL_X32 FILLER_0_56_1108 ();
 FILLCELL_X8 FILLER_0_56_1140 ();
 FILLCELL_X32 FILLER_0_57_1 ();
 FILLCELL_X32 FILLER_0_57_33 ();
 FILLCELL_X32 FILLER_0_57_65 ();
 FILLCELL_X32 FILLER_0_57_97 ();
 FILLCELL_X16 FILLER_0_57_129 ();
 FILLCELL_X8 FILLER_0_57_145 ();
 FILLCELL_X4 FILLER_0_57_153 ();
 FILLCELL_X1 FILLER_0_57_216 ();
 FILLCELL_X2 FILLER_0_57_234 ();
 FILLCELL_X1 FILLER_0_57_246 ();
 FILLCELL_X1 FILLER_0_57_335 ();
 FILLCELL_X1 FILLER_0_57_353 ();
 FILLCELL_X2 FILLER_0_57_364 ();
 FILLCELL_X1 FILLER_0_57_366 ();
 FILLCELL_X1 FILLER_0_57_407 ();
 FILLCELL_X1 FILLER_0_57_417 ();
 FILLCELL_X2 FILLER_0_57_440 ();
 FILLCELL_X1 FILLER_0_57_457 ();
 FILLCELL_X1 FILLER_0_57_463 ();
 FILLCELL_X4 FILLER_0_57_474 ();
 FILLCELL_X2 FILLER_0_57_497 ();
 FILLCELL_X1 FILLER_0_57_499 ();
 FILLCELL_X1 FILLER_0_57_517 ();
 FILLCELL_X1 FILLER_0_57_543 ();
 FILLCELL_X1 FILLER_0_57_564 ();
 FILLCELL_X1 FILLER_0_57_570 ();
 FILLCELL_X2 FILLER_0_57_604 ();
 FILLCELL_X1 FILLER_0_57_606 ();
 FILLCELL_X1 FILLER_0_57_634 ();
 FILLCELL_X2 FILLER_0_57_645 ();
 FILLCELL_X8 FILLER_0_57_670 ();
 FILLCELL_X2 FILLER_0_57_678 ();
 FILLCELL_X1 FILLER_0_57_680 ();
 FILLCELL_X4 FILLER_0_57_716 ();
 FILLCELL_X4 FILLER_0_57_724 ();
 FILLCELL_X1 FILLER_0_57_728 ();
 FILLCELL_X8 FILLER_0_57_749 ();
 FILLCELL_X4 FILLER_0_57_757 ();
 FILLCELL_X2 FILLER_0_57_771 ();
 FILLCELL_X1 FILLER_0_57_773 ();
 FILLCELL_X1 FILLER_0_57_807 ();
 FILLCELL_X4 FILLER_0_57_832 ();
 FILLCELL_X2 FILLER_0_57_842 ();
 FILLCELL_X1 FILLER_0_57_844 ();
 FILLCELL_X1 FILLER_0_57_859 ();
 FILLCELL_X2 FILLER_0_57_874 ();
 FILLCELL_X1 FILLER_0_57_891 ();
 FILLCELL_X1 FILLER_0_57_902 ();
 FILLCELL_X2 FILLER_0_57_908 ();
 FILLCELL_X2 FILLER_0_57_917 ();
 FILLCELL_X2 FILLER_0_57_935 ();
 FILLCELL_X1 FILLER_0_57_954 ();
 FILLCELL_X4 FILLER_0_57_972 ();
 FILLCELL_X1 FILLER_0_57_999 ();
 FILLCELL_X1 FILLER_0_57_1010 ();
 FILLCELL_X1 FILLER_0_57_1016 ();
 FILLCELL_X1 FILLER_0_57_1027 ();
 FILLCELL_X1 FILLER_0_57_1038 ();
 FILLCELL_X1 FILLER_0_57_1049 ();
 FILLCELL_X32 FILLER_0_57_1079 ();
 FILLCELL_X32 FILLER_0_57_1111 ();
 FILLCELL_X4 FILLER_0_57_1143 ();
 FILLCELL_X1 FILLER_0_57_1147 ();
 FILLCELL_X32 FILLER_0_58_1 ();
 FILLCELL_X32 FILLER_0_58_33 ();
 FILLCELL_X32 FILLER_0_58_65 ();
 FILLCELL_X32 FILLER_0_58_97 ();
 FILLCELL_X32 FILLER_0_58_129 ();
 FILLCELL_X8 FILLER_0_58_161 ();
 FILLCELL_X1 FILLER_0_58_169 ();
 FILLCELL_X4 FILLER_0_58_180 ();
 FILLCELL_X4 FILLER_0_58_294 ();
 FILLCELL_X1 FILLER_0_58_318 ();
 FILLCELL_X1 FILLER_0_58_383 ();
 FILLCELL_X1 FILLER_0_58_421 ();
 FILLCELL_X1 FILLER_0_58_426 ();
 FILLCELL_X1 FILLER_0_58_437 ();
 FILLCELL_X4 FILLER_0_58_450 ();
 FILLCELL_X2 FILLER_0_58_454 ();
 FILLCELL_X2 FILLER_0_58_466 ();
 FILLCELL_X1 FILLER_0_58_468 ();
 FILLCELL_X4 FILLER_0_58_474 ();
 FILLCELL_X1 FILLER_0_58_478 ();
 FILLCELL_X2 FILLER_0_58_485 ();
 FILLCELL_X1 FILLER_0_58_538 ();
 FILLCELL_X1 FILLER_0_58_566 ();
 FILLCELL_X2 FILLER_0_58_592 ();
 FILLCELL_X1 FILLER_0_58_604 ();
 FILLCELL_X2 FILLER_0_58_629 ();
 FILLCELL_X1 FILLER_0_58_651 ();
 FILLCELL_X2 FILLER_0_58_675 ();
 FILLCELL_X1 FILLER_0_58_677 ();
 FILLCELL_X4 FILLER_0_58_682 ();
 FILLCELL_X2 FILLER_0_58_686 ();
 FILLCELL_X1 FILLER_0_58_733 ();
 FILLCELL_X1 FILLER_0_58_744 ();
 FILLCELL_X2 FILLER_0_58_761 ();
 FILLCELL_X2 FILLER_0_58_796 ();
 FILLCELL_X4 FILLER_0_58_811 ();
 FILLCELL_X1 FILLER_0_58_815 ();
 FILLCELL_X1 FILLER_0_58_821 ();
 FILLCELL_X1 FILLER_0_58_824 ();
 FILLCELL_X2 FILLER_0_58_849 ();
 FILLCELL_X1 FILLER_0_58_851 ();
 FILLCELL_X2 FILLER_0_58_867 ();
 FILLCELL_X1 FILLER_0_58_869 ();
 FILLCELL_X2 FILLER_0_58_899 ();
 FILLCELL_X1 FILLER_0_58_901 ();
 FILLCELL_X4 FILLER_0_58_926 ();
 FILLCELL_X2 FILLER_0_58_964 ();
 FILLCELL_X2 FILLER_0_58_1003 ();
 FILLCELL_X32 FILLER_0_58_1077 ();
 FILLCELL_X1 FILLER_0_58_1109 ();
 FILLCELL_X16 FILLER_0_58_1120 ();
 FILLCELL_X8 FILLER_0_58_1136 ();
 FILLCELL_X4 FILLER_0_58_1144 ();
 FILLCELL_X32 FILLER_0_59_1 ();
 FILLCELL_X32 FILLER_0_59_33 ();
 FILLCELL_X32 FILLER_0_59_65 ();
 FILLCELL_X32 FILLER_0_59_97 ();
 FILLCELL_X16 FILLER_0_59_129 ();
 FILLCELL_X8 FILLER_0_59_145 ();
 FILLCELL_X2 FILLER_0_59_153 ();
 FILLCELL_X1 FILLER_0_59_155 ();
 FILLCELL_X8 FILLER_0_59_166 ();
 FILLCELL_X4 FILLER_0_59_174 ();
 FILLCELL_X2 FILLER_0_59_178 ();
 FILLCELL_X2 FILLER_0_59_199 ();
 FILLCELL_X1 FILLER_0_59_218 ();
 FILLCELL_X1 FILLER_0_59_257 ();
 FILLCELL_X2 FILLER_0_59_285 ();
 FILLCELL_X1 FILLER_0_59_287 ();
 FILLCELL_X2 FILLER_0_59_319 ();
 FILLCELL_X2 FILLER_0_59_355 ();
 FILLCELL_X2 FILLER_0_59_388 ();
 FILLCELL_X2 FILLER_0_59_400 ();
 FILLCELL_X1 FILLER_0_59_434 ();
 FILLCELL_X2 FILLER_0_59_458 ();
 FILLCELL_X8 FILLER_0_59_482 ();
 FILLCELL_X1 FILLER_0_59_503 ();
 FILLCELL_X1 FILLER_0_59_514 ();
 FILLCELL_X1 FILLER_0_59_536 ();
 FILLCELL_X1 FILLER_0_59_559 ();
 FILLCELL_X1 FILLER_0_59_579 ();
 FILLCELL_X2 FILLER_0_59_611 ();
 FILLCELL_X1 FILLER_0_59_689 ();
 FILLCELL_X2 FILLER_0_59_712 ();
 FILLCELL_X1 FILLER_0_59_714 ();
 FILLCELL_X2 FILLER_0_59_729 ();
 FILLCELL_X4 FILLER_0_59_739 ();
 FILLCELL_X2 FILLER_0_59_743 ();
 FILLCELL_X1 FILLER_0_59_745 ();
 FILLCELL_X1 FILLER_0_59_761 ();
 FILLCELL_X1 FILLER_0_59_791 ();
 FILLCELL_X4 FILLER_0_59_811 ();
 FILLCELL_X1 FILLER_0_59_815 ();
 FILLCELL_X2 FILLER_0_59_828 ();
 FILLCELL_X1 FILLER_0_59_830 ();
 FILLCELL_X1 FILLER_0_59_848 ();
 FILLCELL_X1 FILLER_0_59_885 ();
 FILLCELL_X2 FILLER_0_59_918 ();
 FILLCELL_X1 FILLER_0_59_940 ();
 FILLCELL_X2 FILLER_0_59_955 ();
 FILLCELL_X4 FILLER_0_59_966 ();
 FILLCELL_X1 FILLER_0_59_977 ();
 FILLCELL_X2 FILLER_0_59_998 ();
 FILLCELL_X1 FILLER_0_59_1010 ();
 FILLCELL_X1 FILLER_0_59_1021 ();
 FILLCELL_X1 FILLER_0_59_1031 ();
 FILLCELL_X2 FILLER_0_59_1037 ();
 FILLCELL_X1 FILLER_0_59_1049 ();
 FILLCELL_X2 FILLER_0_59_1059 ();
 FILLCELL_X1 FILLER_0_59_1061 ();
 FILLCELL_X4 FILLER_0_59_1067 ();
 FILLCELL_X16 FILLER_0_59_1081 ();
 FILLCELL_X4 FILLER_0_59_1097 ();
 FILLCELL_X1 FILLER_0_59_1101 ();
 FILLCELL_X8 FILLER_0_59_1138 ();
 FILLCELL_X2 FILLER_0_59_1146 ();
 FILLCELL_X32 FILLER_0_60_1 ();
 FILLCELL_X32 FILLER_0_60_33 ();
 FILLCELL_X32 FILLER_0_60_65 ();
 FILLCELL_X32 FILLER_0_60_97 ();
 FILLCELL_X16 FILLER_0_60_129 ();
 FILLCELL_X8 FILLER_0_60_145 ();
 FILLCELL_X4 FILLER_0_60_153 ();
 FILLCELL_X1 FILLER_0_60_196 ();
 FILLCELL_X1 FILLER_0_60_219 ();
 FILLCELL_X2 FILLER_0_60_239 ();
 FILLCELL_X1 FILLER_0_60_251 ();
 FILLCELL_X1 FILLER_0_60_276 ();
 FILLCELL_X1 FILLER_0_60_301 ();
 FILLCELL_X1 FILLER_0_60_319 ();
 FILLCELL_X1 FILLER_0_60_355 ();
 FILLCELL_X1 FILLER_0_60_394 ();
 FILLCELL_X2 FILLER_0_60_410 ();
 FILLCELL_X2 FILLER_0_60_427 ();
 FILLCELL_X1 FILLER_0_60_444 ();
 FILLCELL_X2 FILLER_0_60_452 ();
 FILLCELL_X4 FILLER_0_60_471 ();
 FILLCELL_X4 FILLER_0_60_484 ();
 FILLCELL_X2 FILLER_0_60_501 ();
 FILLCELL_X1 FILLER_0_60_517 ();
 FILLCELL_X1 FILLER_0_60_567 ();
 FILLCELL_X2 FILLER_0_60_603 ();
 FILLCELL_X1 FILLER_0_60_656 ();
 FILLCELL_X1 FILLER_0_60_716 ();
 FILLCELL_X2 FILLER_0_60_784 ();
 FILLCELL_X2 FILLER_0_60_791 ();
 FILLCELL_X1 FILLER_0_60_796 ();
 FILLCELL_X1 FILLER_0_60_807 ();
 FILLCELL_X1 FILLER_0_60_812 ();
 FILLCELL_X8 FILLER_0_60_816 ();
 FILLCELL_X1 FILLER_0_60_834 ();
 FILLCELL_X1 FILLER_0_60_856 ();
 FILLCELL_X1 FILLER_0_60_909 ();
 FILLCELL_X4 FILLER_0_60_920 ();
 FILLCELL_X2 FILLER_0_60_924 ();
 FILLCELL_X1 FILLER_0_60_926 ();
 FILLCELL_X2 FILLER_0_60_962 ();
 FILLCELL_X2 FILLER_0_60_974 ();
 FILLCELL_X1 FILLER_0_60_976 ();
 FILLCELL_X2 FILLER_0_60_1026 ();
 FILLCELL_X8 FILLER_0_60_1038 ();
 FILLCELL_X8 FILLER_0_60_1071 ();
 FILLCELL_X4 FILLER_0_60_1099 ();
 FILLCELL_X1 FILLER_0_60_1103 ();
 FILLCELL_X32 FILLER_0_61_1 ();
 FILLCELL_X32 FILLER_0_61_33 ();
 FILLCELL_X32 FILLER_0_61_65 ();
 FILLCELL_X32 FILLER_0_61_97 ();
 FILLCELL_X32 FILLER_0_61_129 ();
 FILLCELL_X1 FILLER_0_61_161 ();
 FILLCELL_X4 FILLER_0_61_232 ();
 FILLCELL_X1 FILLER_0_61_246 ();
 FILLCELL_X1 FILLER_0_61_262 ();
 FILLCELL_X1 FILLER_0_61_273 ();
 FILLCELL_X1 FILLER_0_61_308 ();
 FILLCELL_X2 FILLER_0_61_350 ();
 FILLCELL_X1 FILLER_0_61_352 ();
 FILLCELL_X2 FILLER_0_61_384 ();
 FILLCELL_X2 FILLER_0_61_409 ();
 FILLCELL_X1 FILLER_0_61_421 ();
 FILLCELL_X1 FILLER_0_61_427 ();
 FILLCELL_X4 FILLER_0_61_438 ();
 FILLCELL_X2 FILLER_0_61_442 ();
 FILLCELL_X1 FILLER_0_61_444 ();
 FILLCELL_X1 FILLER_0_61_486 ();
 FILLCELL_X1 FILLER_0_61_556 ();
 FILLCELL_X1 FILLER_0_61_592 ();
 FILLCELL_X1 FILLER_0_61_622 ();
 FILLCELL_X1 FILLER_0_61_681 ();
 FILLCELL_X2 FILLER_0_61_696 ();
 FILLCELL_X1 FILLER_0_61_727 ();
 FILLCELL_X1 FILLER_0_61_732 ();
 FILLCELL_X1 FILLER_0_61_748 ();
 FILLCELL_X2 FILLER_0_61_784 ();
 FILLCELL_X8 FILLER_0_61_796 ();
 FILLCELL_X1 FILLER_0_61_835 ();
 FILLCELL_X2 FILLER_0_61_851 ();
 FILLCELL_X8 FILLER_0_61_920 ();
 FILLCELL_X1 FILLER_0_61_928 ();
 FILLCELL_X4 FILLER_0_61_971 ();
 FILLCELL_X1 FILLER_0_61_985 ();
 FILLCELL_X8 FILLER_0_61_1005 ();
 FILLCELL_X1 FILLER_0_61_1023 ();
 FILLCELL_X2 FILLER_0_61_1029 ();
 FILLCELL_X1 FILLER_0_61_1031 ();
 FILLCELL_X16 FILLER_0_61_1052 ();
 FILLCELL_X4 FILLER_0_61_1068 ();
 FILLCELL_X1 FILLER_0_61_1072 ();
 FILLCELL_X1 FILLER_0_61_1096 ();
 FILLCELL_X1 FILLER_0_61_1120 ();
 FILLCELL_X8 FILLER_0_61_1140 ();
 FILLCELL_X32 FILLER_0_62_1 ();
 FILLCELL_X32 FILLER_0_62_33 ();
 FILLCELL_X32 FILLER_0_62_65 ();
 FILLCELL_X32 FILLER_0_62_97 ();
 FILLCELL_X32 FILLER_0_62_129 ();
 FILLCELL_X4 FILLER_0_62_161 ();
 FILLCELL_X1 FILLER_0_62_165 ();
 FILLCELL_X1 FILLER_0_62_176 ();
 FILLCELL_X2 FILLER_0_62_202 ();
 FILLCELL_X1 FILLER_0_62_204 ();
 FILLCELL_X4 FILLER_0_62_215 ();
 FILLCELL_X2 FILLER_0_62_224 ();
 FILLCELL_X1 FILLER_0_62_271 ();
 FILLCELL_X1 FILLER_0_62_299 ();
 FILLCELL_X4 FILLER_0_62_390 ();
 FILLCELL_X2 FILLER_0_62_408 ();
 FILLCELL_X2 FILLER_0_62_414 ();
 FILLCELL_X4 FILLER_0_62_436 ();
 FILLCELL_X2 FILLER_0_62_483 ();
 FILLCELL_X1 FILLER_0_62_520 ();
 FILLCELL_X1 FILLER_0_62_528 ();
 FILLCELL_X2 FILLER_0_62_606 ();
 FILLCELL_X2 FILLER_0_62_629 ();
 FILLCELL_X2 FILLER_0_62_639 ();
 FILLCELL_X1 FILLER_0_62_641 ();
 FILLCELL_X2 FILLER_0_62_669 ();
 FILLCELL_X1 FILLER_0_62_694 ();
 FILLCELL_X2 FILLER_0_62_742 ();
 FILLCELL_X2 FILLER_0_62_753 ();
 FILLCELL_X1 FILLER_0_62_773 ();
 FILLCELL_X8 FILLER_0_62_805 ();
 FILLCELL_X4 FILLER_0_62_813 ();
 FILLCELL_X1 FILLER_0_62_817 ();
 FILLCELL_X2 FILLER_0_62_841 ();
 FILLCELL_X2 FILLER_0_62_894 ();
 FILLCELL_X4 FILLER_0_62_906 ();
 FILLCELL_X2 FILLER_0_62_937 ();
 FILLCELL_X1 FILLER_0_62_939 ();
 FILLCELL_X2 FILLER_0_62_945 ();
 FILLCELL_X1 FILLER_0_62_947 ();
 FILLCELL_X8 FILLER_0_62_968 ();
 FILLCELL_X4 FILLER_0_62_976 ();
 FILLCELL_X1 FILLER_0_62_980 ();
 FILLCELL_X16 FILLER_0_62_1001 ();
 FILLCELL_X2 FILLER_0_62_1017 ();
 FILLCELL_X4 FILLER_0_62_1029 ();
 FILLCELL_X1 FILLER_0_62_1033 ();
 FILLCELL_X2 FILLER_0_62_1039 ();
 FILLCELL_X8 FILLER_0_62_1051 ();
 FILLCELL_X4 FILLER_0_62_1059 ();
 FILLCELL_X2 FILLER_0_62_1063 ();
 FILLCELL_X1 FILLER_0_62_1065 ();
 FILLCELL_X1 FILLER_0_62_1102 ();
 FILLCELL_X1 FILLER_0_62_1107 ();
 FILLCELL_X1 FILLER_0_62_1112 ();
 FILLCELL_X1 FILLER_0_62_1116 ();
 FILLCELL_X1 FILLER_0_62_1122 ();
 FILLCELL_X1 FILLER_0_62_1132 ();
 FILLCELL_X1 FILLER_0_62_1137 ();
 FILLCELL_X32 FILLER_0_63_1 ();
 FILLCELL_X32 FILLER_0_63_33 ();
 FILLCELL_X32 FILLER_0_63_65 ();
 FILLCELL_X32 FILLER_0_63_97 ();
 FILLCELL_X32 FILLER_0_63_129 ();
 FILLCELL_X4 FILLER_0_63_161 ();
 FILLCELL_X2 FILLER_0_63_165 ();
 FILLCELL_X1 FILLER_0_63_167 ();
 FILLCELL_X8 FILLER_0_63_178 ();
 FILLCELL_X4 FILLER_0_63_186 ();
 FILLCELL_X2 FILLER_0_63_190 ();
 FILLCELL_X4 FILLER_0_63_202 ();
 FILLCELL_X2 FILLER_0_63_211 ();
 FILLCELL_X2 FILLER_0_63_254 ();
 FILLCELL_X2 FILLER_0_63_266 ();
 FILLCELL_X2 FILLER_0_63_278 ();
 FILLCELL_X1 FILLER_0_63_280 ();
 FILLCELL_X2 FILLER_0_63_302 ();
 FILLCELL_X2 FILLER_0_63_319 ();
 FILLCELL_X2 FILLER_0_63_355 ();
 FILLCELL_X2 FILLER_0_63_364 ();
 FILLCELL_X1 FILLER_0_63_400 ();
 FILLCELL_X1 FILLER_0_63_423 ();
 FILLCELL_X2 FILLER_0_63_434 ();
 FILLCELL_X1 FILLER_0_63_436 ();
 FILLCELL_X1 FILLER_0_63_603 ();
 FILLCELL_X1 FILLER_0_63_614 ();
 FILLCELL_X1 FILLER_0_63_677 ();
 FILLCELL_X1 FILLER_0_63_688 ();
 FILLCELL_X1 FILLER_0_63_726 ();
 FILLCELL_X1 FILLER_0_63_731 ();
 FILLCELL_X1 FILLER_0_63_737 ();
 FILLCELL_X2 FILLER_0_63_747 ();
 FILLCELL_X2 FILLER_0_63_793 ();
 FILLCELL_X2 FILLER_0_63_815 ();
 FILLCELL_X1 FILLER_0_63_861 ();
 FILLCELL_X2 FILLER_0_63_867 ();
 FILLCELL_X2 FILLER_0_63_928 ();
 FILLCELL_X1 FILLER_0_63_930 ();
 FILLCELL_X8 FILLER_0_63_941 ();
 FILLCELL_X1 FILLER_0_63_949 ();
 FILLCELL_X2 FILLER_0_63_955 ();
 FILLCELL_X2 FILLER_0_63_967 ();
 FILLCELL_X4 FILLER_0_63_979 ();
 FILLCELL_X2 FILLER_0_63_983 ();
 FILLCELL_X1 FILLER_0_63_1009 ();
 FILLCELL_X4 FILLER_0_63_1015 ();
 FILLCELL_X1 FILLER_0_63_1019 ();
 FILLCELL_X32 FILLER_0_63_1045 ();
 FILLCELL_X1 FILLER_0_63_1077 ();
 FILLCELL_X2 FILLER_0_63_1111 ();
 FILLCELL_X8 FILLER_0_63_1137 ();
 FILLCELL_X2 FILLER_0_63_1145 ();
 FILLCELL_X1 FILLER_0_63_1147 ();
 FILLCELL_X32 FILLER_0_64_1 ();
 FILLCELL_X32 FILLER_0_64_33 ();
 FILLCELL_X32 FILLER_0_64_65 ();
 FILLCELL_X32 FILLER_0_64_97 ();
 FILLCELL_X32 FILLER_0_64_129 ();
 FILLCELL_X1 FILLER_0_64_161 ();
 FILLCELL_X1 FILLER_0_64_177 ();
 FILLCELL_X8 FILLER_0_64_187 ();
 FILLCELL_X1 FILLER_0_64_195 ();
 FILLCELL_X8 FILLER_0_64_206 ();
 FILLCELL_X2 FILLER_0_64_214 ();
 FILLCELL_X1 FILLER_0_64_216 ();
 FILLCELL_X8 FILLER_0_64_222 ();
 FILLCELL_X1 FILLER_0_64_230 ();
 FILLCELL_X2 FILLER_0_64_241 ();
 FILLCELL_X2 FILLER_0_64_347 ();
 FILLCELL_X2 FILLER_0_64_359 ();
 FILLCELL_X1 FILLER_0_64_361 ();
 FILLCELL_X2 FILLER_0_64_369 ();
 FILLCELL_X2 FILLER_0_64_377 ();
 FILLCELL_X2 FILLER_0_64_384 ();
 FILLCELL_X2 FILLER_0_64_425 ();
 FILLCELL_X4 FILLER_0_64_435 ();
 FILLCELL_X1 FILLER_0_64_439 ();
 FILLCELL_X8 FILLER_0_64_443 ();
 FILLCELL_X1 FILLER_0_64_451 ();
 FILLCELL_X2 FILLER_0_64_617 ();
 FILLCELL_X1 FILLER_0_64_619 ();
 FILLCELL_X1 FILLER_0_64_630 ();
 FILLCELL_X2 FILLER_0_64_646 ();
 FILLCELL_X1 FILLER_0_64_648 ();
 FILLCELL_X1 FILLER_0_64_681 ();
 FILLCELL_X2 FILLER_0_64_699 ();
 FILLCELL_X2 FILLER_0_64_720 ();
 FILLCELL_X4 FILLER_0_64_725 ();
 FILLCELL_X1 FILLER_0_64_793 ();
 FILLCELL_X2 FILLER_0_64_824 ();
 FILLCELL_X2 FILLER_0_64_877 ();
 FILLCELL_X1 FILLER_0_64_904 ();
 FILLCELL_X1 FILLER_0_64_930 ();
 FILLCELL_X2 FILLER_0_64_941 ();
 FILLCELL_X2 FILLER_0_64_948 ();
 FILLCELL_X1 FILLER_0_64_960 ();
 FILLCELL_X1 FILLER_0_64_978 ();
 FILLCELL_X1 FILLER_0_64_994 ();
 FILLCELL_X1 FILLER_0_64_1005 ();
 FILLCELL_X1 FILLER_0_64_1016 ();
 FILLCELL_X16 FILLER_0_64_1027 ();
 FILLCELL_X8 FILLER_0_64_1043 ();
 FILLCELL_X4 FILLER_0_64_1051 ();
 FILLCELL_X1 FILLER_0_64_1055 ();
 FILLCELL_X16 FILLER_0_64_1076 ();
 FILLCELL_X8 FILLER_0_64_1092 ();
 FILLCELL_X2 FILLER_0_64_1100 ();
 FILLCELL_X1 FILLER_0_64_1109 ();
 FILLCELL_X2 FILLER_0_64_1126 ();
 FILLCELL_X32 FILLER_0_65_1 ();
 FILLCELL_X32 FILLER_0_65_33 ();
 FILLCELL_X32 FILLER_0_65_65 ();
 FILLCELL_X32 FILLER_0_65_97 ();
 FILLCELL_X32 FILLER_0_65_129 ();
 FILLCELL_X1 FILLER_0_65_161 ();
 FILLCELL_X1 FILLER_0_65_172 ();
 FILLCELL_X2 FILLER_0_65_178 ();
 FILLCELL_X1 FILLER_0_65_190 ();
 FILLCELL_X2 FILLER_0_65_200 ();
 FILLCELL_X1 FILLER_0_65_202 ();
 FILLCELL_X1 FILLER_0_65_213 ();
 FILLCELL_X4 FILLER_0_65_224 ();
 FILLCELL_X2 FILLER_0_65_247 ();
 FILLCELL_X1 FILLER_0_65_249 ();
 FILLCELL_X2 FILLER_0_65_260 ();
 FILLCELL_X1 FILLER_0_65_262 ();
 FILLCELL_X2 FILLER_0_65_278 ();
 FILLCELL_X1 FILLER_0_65_280 ();
 FILLCELL_X4 FILLER_0_65_286 ();
 FILLCELL_X2 FILLER_0_65_305 ();
 FILLCELL_X1 FILLER_0_65_307 ();
 FILLCELL_X2 FILLER_0_65_390 ();
 FILLCELL_X1 FILLER_0_65_392 ();
 FILLCELL_X2 FILLER_0_65_413 ();
 FILLCELL_X1 FILLER_0_65_425 ();
 FILLCELL_X2 FILLER_0_65_440 ();
 FILLCELL_X1 FILLER_0_65_449 ();
 FILLCELL_X2 FILLER_0_65_477 ();
 FILLCELL_X1 FILLER_0_65_598 ();
 FILLCELL_X1 FILLER_0_65_655 ();
 FILLCELL_X1 FILLER_0_65_680 ();
 FILLCELL_X1 FILLER_0_65_696 ();
 FILLCELL_X1 FILLER_0_65_744 ();
 FILLCELL_X1 FILLER_0_65_792 ();
 FILLCELL_X4 FILLER_0_65_813 ();
 FILLCELL_X1 FILLER_0_65_817 ();
 FILLCELL_X2 FILLER_0_65_822 ();
 FILLCELL_X1 FILLER_0_65_833 ();
 FILLCELL_X2 FILLER_0_65_844 ();
 FILLCELL_X2 FILLER_0_65_856 ();
 FILLCELL_X1 FILLER_0_65_865 ();
 FILLCELL_X2 FILLER_0_65_923 ();
 FILLCELL_X8 FILLER_0_65_935 ();
 FILLCELL_X2 FILLER_0_65_943 ();
 FILLCELL_X4 FILLER_0_65_960 ();
 FILLCELL_X4 FILLER_0_65_974 ();
 FILLCELL_X2 FILLER_0_65_978 ();
 FILLCELL_X4 FILLER_0_65_990 ();
 FILLCELL_X2 FILLER_0_65_994 ();
 FILLCELL_X1 FILLER_0_65_996 ();
 FILLCELL_X16 FILLER_0_65_1017 ();
 FILLCELL_X4 FILLER_0_65_1033 ();
 FILLCELL_X1 FILLER_0_65_1059 ();
 FILLCELL_X1 FILLER_0_65_1103 ();
 FILLCELL_X2 FILLER_0_65_1124 ();
 FILLCELL_X2 FILLER_0_65_1146 ();
 FILLCELL_X32 FILLER_0_66_1 ();
 FILLCELL_X32 FILLER_0_66_33 ();
 FILLCELL_X32 FILLER_0_66_65 ();
 FILLCELL_X32 FILLER_0_66_97 ();
 FILLCELL_X32 FILLER_0_66_129 ();
 FILLCELL_X2 FILLER_0_66_201 ();
 FILLCELL_X1 FILLER_0_66_203 ();
 FILLCELL_X2 FILLER_0_66_233 ();
 FILLCELL_X1 FILLER_0_66_265 ();
 FILLCELL_X4 FILLER_0_66_291 ();
 FILLCELL_X1 FILLER_0_66_295 ();
 FILLCELL_X2 FILLER_0_66_305 ();
 FILLCELL_X8 FILLER_0_66_342 ();
 FILLCELL_X1 FILLER_0_66_350 ();
 FILLCELL_X1 FILLER_0_66_382 ();
 FILLCELL_X4 FILLER_0_66_393 ();
 FILLCELL_X8 FILLER_0_66_400 ();
 FILLCELL_X1 FILLER_0_66_408 ();
 FILLCELL_X1 FILLER_0_66_460 ();
 FILLCELL_X1 FILLER_0_66_471 ();
 FILLCELL_X1 FILLER_0_66_513 ();
 FILLCELL_X1 FILLER_0_66_546 ();
 FILLCELL_X1 FILLER_0_66_594 ();
 FILLCELL_X1 FILLER_0_66_630 ();
 FILLCELL_X1 FILLER_0_66_685 ();
 FILLCELL_X2 FILLER_0_66_708 ();
 FILLCELL_X1 FILLER_0_66_729 ();
 FILLCELL_X1 FILLER_0_66_786 ();
 FILLCELL_X1 FILLER_0_66_793 ();
 FILLCELL_X2 FILLER_0_66_814 ();
 FILLCELL_X1 FILLER_0_66_816 ();
 FILLCELL_X2 FILLER_0_66_869 ();
 FILLCELL_X8 FILLER_0_66_912 ();
 FILLCELL_X32 FILLER_0_66_925 ();
 FILLCELL_X16 FILLER_0_66_957 ();
 FILLCELL_X4 FILLER_0_66_973 ();
 FILLCELL_X2 FILLER_0_66_977 ();
 FILLCELL_X4 FILLER_0_66_984 ();
 FILLCELL_X1 FILLER_0_66_988 ();
 FILLCELL_X2 FILLER_0_66_1008 ();
 FILLCELL_X1 FILLER_0_66_1010 ();
 FILLCELL_X1 FILLER_0_66_1016 ();
 FILLCELL_X4 FILLER_0_66_1027 ();
 FILLCELL_X2 FILLER_0_66_1031 ();
 FILLCELL_X1 FILLER_0_66_1033 ();
 FILLCELL_X4 FILLER_0_66_1116 ();
 FILLCELL_X4 FILLER_0_66_1141 ();
 FILLCELL_X2 FILLER_0_66_1145 ();
 FILLCELL_X1 FILLER_0_66_1147 ();
 FILLCELL_X32 FILLER_0_67_1 ();
 FILLCELL_X32 FILLER_0_67_33 ();
 FILLCELL_X32 FILLER_0_67_65 ();
 FILLCELL_X32 FILLER_0_67_97 ();
 FILLCELL_X32 FILLER_0_67_129 ();
 FILLCELL_X4 FILLER_0_67_161 ();
 FILLCELL_X4 FILLER_0_67_185 ();
 FILLCELL_X1 FILLER_0_67_199 ();
 FILLCELL_X2 FILLER_0_67_205 ();
 FILLCELL_X1 FILLER_0_67_207 ();
 FILLCELL_X2 FILLER_0_67_218 ();
 FILLCELL_X1 FILLER_0_67_220 ();
 FILLCELL_X1 FILLER_0_67_240 ();
 FILLCELL_X1 FILLER_0_67_260 ();
 FILLCELL_X16 FILLER_0_67_286 ();
 FILLCELL_X2 FILLER_0_67_302 ();
 FILLCELL_X8 FILLER_0_67_337 ();
 FILLCELL_X4 FILLER_0_67_345 ();
 FILLCELL_X2 FILLER_0_67_362 ();
 FILLCELL_X1 FILLER_0_67_369 ();
 FILLCELL_X8 FILLER_0_67_380 ();
 FILLCELL_X4 FILLER_0_67_388 ();
 FILLCELL_X1 FILLER_0_67_392 ();
 FILLCELL_X2 FILLER_0_67_435 ();
 FILLCELL_X2 FILLER_0_67_509 ();
 FILLCELL_X1 FILLER_0_67_511 ();
 FILLCELL_X2 FILLER_0_67_530 ();
 FILLCELL_X2 FILLER_0_67_659 ();
 FILLCELL_X1 FILLER_0_67_661 ();
 FILLCELL_X2 FILLER_0_67_672 ();
 FILLCELL_X1 FILLER_0_67_674 ();
 FILLCELL_X1 FILLER_0_67_716 ();
 FILLCELL_X1 FILLER_0_67_763 ();
 FILLCELL_X8 FILLER_0_67_807 ();
 FILLCELL_X4 FILLER_0_67_815 ();
 FILLCELL_X1 FILLER_0_67_826 ();
 FILLCELL_X2 FILLER_0_67_834 ();
 FILLCELL_X1 FILLER_0_67_847 ();
 FILLCELL_X1 FILLER_0_67_855 ();
 FILLCELL_X1 FILLER_0_67_886 ();
 FILLCELL_X1 FILLER_0_67_909 ();
 FILLCELL_X4 FILLER_0_67_932 ();
 FILLCELL_X4 FILLER_0_67_941 ();
 FILLCELL_X2 FILLER_0_67_945 ();
 FILLCELL_X2 FILLER_0_67_952 ();
 FILLCELL_X2 FILLER_0_67_978 ();
 FILLCELL_X16 FILLER_0_67_1039 ();
 FILLCELL_X8 FILLER_0_67_1110 ();
 FILLCELL_X2 FILLER_0_67_1118 ();
 FILLCELL_X1 FILLER_0_67_1120 ();
 FILLCELL_X2 FILLER_0_67_1125 ();
 FILLCELL_X1 FILLER_0_67_1127 ();
 FILLCELL_X8 FILLER_0_67_1135 ();
 FILLCELL_X4 FILLER_0_67_1143 ();
 FILLCELL_X1 FILLER_0_67_1147 ();
 FILLCELL_X32 FILLER_0_68_1 ();
 FILLCELL_X32 FILLER_0_68_33 ();
 FILLCELL_X32 FILLER_0_68_65 ();
 FILLCELL_X32 FILLER_0_68_97 ();
 FILLCELL_X32 FILLER_0_68_129 ();
 FILLCELL_X16 FILLER_0_68_161 ();
 FILLCELL_X4 FILLER_0_68_177 ();
 FILLCELL_X2 FILLER_0_68_181 ();
 FILLCELL_X32 FILLER_0_68_193 ();
 FILLCELL_X16 FILLER_0_68_225 ();
 FILLCELL_X4 FILLER_0_68_241 ();
 FILLCELL_X2 FILLER_0_68_255 ();
 FILLCELL_X16 FILLER_0_68_262 ();
 FILLCELL_X4 FILLER_0_68_278 ();
 FILLCELL_X2 FILLER_0_68_282 ();
 FILLCELL_X4 FILLER_0_68_291 ();
 FILLCELL_X2 FILLER_0_68_295 ();
 FILLCELL_X1 FILLER_0_68_297 ();
 FILLCELL_X8 FILLER_0_68_313 ();
 FILLCELL_X2 FILLER_0_68_340 ();
 FILLCELL_X1 FILLER_0_68_342 ();
 FILLCELL_X2 FILLER_0_68_346 ();
 FILLCELL_X4 FILLER_0_68_352 ();
 FILLCELL_X1 FILLER_0_68_356 ();
 FILLCELL_X1 FILLER_0_68_368 ();
 FILLCELL_X16 FILLER_0_68_372 ();
 FILLCELL_X4 FILLER_0_68_388 ();
 FILLCELL_X2 FILLER_0_68_392 ();
 FILLCELL_X2 FILLER_0_68_407 ();
 FILLCELL_X1 FILLER_0_68_420 ();
 FILLCELL_X4 FILLER_0_68_428 ();
 FILLCELL_X1 FILLER_0_68_432 ();
 FILLCELL_X2 FILLER_0_68_443 ();
 FILLCELL_X1 FILLER_0_68_445 ();
 FILLCELL_X1 FILLER_0_68_460 ();
 FILLCELL_X1 FILLER_0_68_491 ();
 FILLCELL_X1 FILLER_0_68_502 ();
 FILLCELL_X2 FILLER_0_68_522 ();
 FILLCELL_X1 FILLER_0_68_534 ();
 FILLCELL_X2 FILLER_0_68_629 ();
 FILLCELL_X1 FILLER_0_68_738 ();
 FILLCELL_X2 FILLER_0_68_786 ();
 FILLCELL_X1 FILLER_0_68_802 ();
 FILLCELL_X4 FILLER_0_68_821 ();
 FILLCELL_X1 FILLER_0_68_835 ();
 FILLCELL_X2 FILLER_0_68_843 ();
 FILLCELL_X2 FILLER_0_68_869 ();
 FILLCELL_X1 FILLER_0_68_924 ();
 FILLCELL_X1 FILLER_0_68_940 ();
 FILLCELL_X2 FILLER_0_68_971 ();
 FILLCELL_X1 FILLER_0_68_973 ();
 FILLCELL_X2 FILLER_0_68_991 ();
 FILLCELL_X8 FILLER_0_68_1030 ();
 FILLCELL_X4 FILLER_0_68_1038 ();
 FILLCELL_X2 FILLER_0_68_1042 ();
 FILLCELL_X1 FILLER_0_68_1075 ();
 FILLCELL_X8 FILLER_0_68_1094 ();
 FILLCELL_X4 FILLER_0_68_1102 ();
 FILLCELL_X2 FILLER_0_68_1106 ();
 FILLCELL_X4 FILLER_0_68_1115 ();
 FILLCELL_X2 FILLER_0_68_1146 ();
 FILLCELL_X32 FILLER_0_69_1 ();
 FILLCELL_X32 FILLER_0_69_33 ();
 FILLCELL_X32 FILLER_0_69_65 ();
 FILLCELL_X32 FILLER_0_69_97 ();
 FILLCELL_X32 FILLER_0_69_129 ();
 FILLCELL_X16 FILLER_0_69_161 ();
 FILLCELL_X8 FILLER_0_69_177 ();
 FILLCELL_X2 FILLER_0_69_194 ();
 FILLCELL_X1 FILLER_0_69_196 ();
 FILLCELL_X16 FILLER_0_69_207 ();
 FILLCELL_X8 FILLER_0_69_223 ();
 FILLCELL_X4 FILLER_0_69_231 ();
 FILLCELL_X4 FILLER_0_69_240 ();
 FILLCELL_X2 FILLER_0_69_244 ();
 FILLCELL_X2 FILLER_0_69_251 ();
 FILLCELL_X2 FILLER_0_69_263 ();
 FILLCELL_X4 FILLER_0_69_270 ();
 FILLCELL_X2 FILLER_0_69_274 ();
 FILLCELL_X1 FILLER_0_69_276 ();
 FILLCELL_X2 FILLER_0_69_350 ();
 FILLCELL_X1 FILLER_0_69_410 ();
 FILLCELL_X1 FILLER_0_69_421 ();
 FILLCELL_X1 FILLER_0_69_432 ();
 FILLCELL_X1 FILLER_0_69_438 ();
 FILLCELL_X1 FILLER_0_69_469 ();
 FILLCELL_X1 FILLER_0_69_486 ();
 FILLCELL_X2 FILLER_0_69_523 ();
 FILLCELL_X4 FILLER_0_69_605 ();
 FILLCELL_X1 FILLER_0_69_636 ();
 FILLCELL_X2 FILLER_0_69_647 ();
 FILLCELL_X1 FILLER_0_69_699 ();
 FILLCELL_X2 FILLER_0_69_710 ();
 FILLCELL_X1 FILLER_0_69_732 ();
 FILLCELL_X2 FILLER_0_69_758 ();
 FILLCELL_X1 FILLER_0_69_760 ();
 FILLCELL_X2 FILLER_0_69_793 ();
 FILLCELL_X1 FILLER_0_69_795 ();
 FILLCELL_X1 FILLER_0_69_809 ();
 FILLCELL_X1 FILLER_0_69_830 ();
 FILLCELL_X1 FILLER_0_69_848 ();
 FILLCELL_X2 FILLER_0_69_856 ();
 FILLCELL_X2 FILLER_0_69_873 ();
 FILLCELL_X1 FILLER_0_69_901 ();
 FILLCELL_X2 FILLER_0_69_924 ();
 FILLCELL_X1 FILLER_0_69_951 ();
 FILLCELL_X1 FILLER_0_69_962 ();
 FILLCELL_X2 FILLER_0_69_973 ();
 FILLCELL_X1 FILLER_0_69_975 ();
 FILLCELL_X4 FILLER_0_69_1010 ();
 FILLCELL_X2 FILLER_0_69_1054 ();
 FILLCELL_X1 FILLER_0_69_1056 ();
 FILLCELL_X1 FILLER_0_69_1086 ();
 FILLCELL_X1 FILLER_0_69_1147 ();
 FILLCELL_X32 FILLER_0_70_1 ();
 FILLCELL_X32 FILLER_0_70_33 ();
 FILLCELL_X32 FILLER_0_70_65 ();
 FILLCELL_X32 FILLER_0_70_97 ();
 FILLCELL_X32 FILLER_0_70_129 ();
 FILLCELL_X8 FILLER_0_70_161 ();
 FILLCELL_X4 FILLER_0_70_169 ();
 FILLCELL_X2 FILLER_0_70_173 ();
 FILLCELL_X2 FILLER_0_70_195 ();
 FILLCELL_X1 FILLER_0_70_202 ();
 FILLCELL_X2 FILLER_0_70_213 ();
 FILLCELL_X2 FILLER_0_70_245 ();
 FILLCELL_X1 FILLER_0_70_294 ();
 FILLCELL_X2 FILLER_0_70_310 ();
 FILLCELL_X2 FILLER_0_70_322 ();
 FILLCELL_X1 FILLER_0_70_334 ();
 FILLCELL_X1 FILLER_0_70_376 ();
 FILLCELL_X1 FILLER_0_70_417 ();
 FILLCELL_X1 FILLER_0_70_462 ();
 FILLCELL_X1 FILLER_0_70_485 ();
 FILLCELL_X1 FILLER_0_70_532 ();
 FILLCELL_X2 FILLER_0_70_654 ();
 FILLCELL_X1 FILLER_0_70_656 ();
 FILLCELL_X4 FILLER_0_70_780 ();
 FILLCELL_X2 FILLER_0_70_784 ();
 FILLCELL_X1 FILLER_0_70_790 ();
 FILLCELL_X2 FILLER_0_70_801 ();
 FILLCELL_X2 FILLER_0_70_825 ();
 FILLCELL_X1 FILLER_0_70_827 ();
 FILLCELL_X4 FILLER_0_70_838 ();
 FILLCELL_X1 FILLER_0_70_842 ();
 FILLCELL_X1 FILLER_0_70_867 ();
 FILLCELL_X1 FILLER_0_70_900 ();
 FILLCELL_X2 FILLER_0_70_938 ();
 FILLCELL_X1 FILLER_0_70_940 ();
 FILLCELL_X1 FILLER_0_70_973 ();
 FILLCELL_X2 FILLER_0_70_983 ();
 FILLCELL_X4 FILLER_0_70_1105 ();
 FILLCELL_X2 FILLER_0_70_1109 ();
 FILLCELL_X1 FILLER_0_70_1121 ();
 FILLCELL_X2 FILLER_0_70_1146 ();
 FILLCELL_X32 FILLER_0_71_1 ();
 FILLCELL_X32 FILLER_0_71_33 ();
 FILLCELL_X32 FILLER_0_71_65 ();
 FILLCELL_X32 FILLER_0_71_97 ();
 FILLCELL_X32 FILLER_0_71_129 ();
 FILLCELL_X8 FILLER_0_71_161 ();
 FILLCELL_X4 FILLER_0_71_169 ();
 FILLCELL_X1 FILLER_0_71_173 ();
 FILLCELL_X8 FILLER_0_71_189 ();
 FILLCELL_X1 FILLER_0_71_206 ();
 FILLCELL_X2 FILLER_0_71_227 ();
 FILLCELL_X1 FILLER_0_71_229 ();
 FILLCELL_X2 FILLER_0_71_245 ();
 FILLCELL_X1 FILLER_0_71_272 ();
 FILLCELL_X2 FILLER_0_71_283 ();
 FILLCELL_X2 FILLER_0_71_319 ();
 FILLCELL_X2 FILLER_0_71_328 ();
 FILLCELL_X2 FILLER_0_71_340 ();
 FILLCELL_X1 FILLER_0_71_384 ();
 FILLCELL_X1 FILLER_0_71_402 ();
 FILLCELL_X1 FILLER_0_71_406 ();
 FILLCELL_X1 FILLER_0_71_417 ();
 FILLCELL_X1 FILLER_0_71_420 ();
 FILLCELL_X1 FILLER_0_71_455 ();
 FILLCELL_X1 FILLER_0_71_505 ();
 FILLCELL_X1 FILLER_0_71_523 ();
 FILLCELL_X1 FILLER_0_71_539 ();
 FILLCELL_X2 FILLER_0_71_569 ();
 FILLCELL_X2 FILLER_0_71_619 ();
 FILLCELL_X2 FILLER_0_71_663 ();
 FILLCELL_X1 FILLER_0_71_713 ();
 FILLCELL_X4 FILLER_0_71_721 ();
 FILLCELL_X1 FILLER_0_71_754 ();
 FILLCELL_X4 FILLER_0_71_799 ();
 FILLCELL_X2 FILLER_0_71_803 ();
 FILLCELL_X1 FILLER_0_71_830 ();
 FILLCELL_X1 FILLER_0_71_845 ();
 FILLCELL_X4 FILLER_0_71_861 ();
 FILLCELL_X2 FILLER_0_71_888 ();
 FILLCELL_X2 FILLER_0_71_900 ();
 FILLCELL_X1 FILLER_0_71_902 ();
 FILLCELL_X2 FILLER_0_71_988 ();
 FILLCELL_X1 FILLER_0_71_990 ();
 FILLCELL_X2 FILLER_0_71_1016 ();
 FILLCELL_X1 FILLER_0_71_1018 ();
 FILLCELL_X1 FILLER_0_71_1080 ();
 FILLCELL_X1 FILLER_0_71_1133 ();
 FILLCELL_X32 FILLER_0_72_1 ();
 FILLCELL_X32 FILLER_0_72_33 ();
 FILLCELL_X32 FILLER_0_72_65 ();
 FILLCELL_X32 FILLER_0_72_97 ();
 FILLCELL_X32 FILLER_0_72_129 ();
 FILLCELL_X16 FILLER_0_72_161 ();
 FILLCELL_X2 FILLER_0_72_177 ();
 FILLCELL_X1 FILLER_0_72_179 ();
 FILLCELL_X2 FILLER_0_72_200 ();
 FILLCELL_X1 FILLER_0_72_202 ();
 FILLCELL_X4 FILLER_0_72_241 ();
 FILLCELL_X1 FILLER_0_72_255 ();
 FILLCELL_X1 FILLER_0_72_290 ();
 FILLCELL_X4 FILLER_0_72_338 ();
 FILLCELL_X2 FILLER_0_72_359 ();
 FILLCELL_X4 FILLER_0_72_439 ();
 FILLCELL_X2 FILLER_0_72_443 ();
 FILLCELL_X4 FILLER_0_72_458 ();
 FILLCELL_X1 FILLER_0_72_462 ();
 FILLCELL_X1 FILLER_0_72_503 ();
 FILLCELL_X2 FILLER_0_72_526 ();
 FILLCELL_X1 FILLER_0_72_572 ();
 FILLCELL_X2 FILLER_0_72_604 ();
 FILLCELL_X1 FILLER_0_72_606 ();
 FILLCELL_X1 FILLER_0_72_681 ();
 FILLCELL_X2 FILLER_0_72_712 ();
 FILLCELL_X2 FILLER_0_72_724 ();
 FILLCELL_X2 FILLER_0_72_753 ();
 FILLCELL_X1 FILLER_0_72_785 ();
 FILLCELL_X8 FILLER_0_72_795 ();
 FILLCELL_X2 FILLER_0_72_803 ();
 FILLCELL_X2 FILLER_0_72_819 ();
 FILLCELL_X2 FILLER_0_72_831 ();
 FILLCELL_X1 FILLER_0_72_843 ();
 FILLCELL_X1 FILLER_0_72_854 ();
 FILLCELL_X2 FILLER_0_72_881 ();
 FILLCELL_X2 FILLER_0_72_922 ();
 FILLCELL_X1 FILLER_0_72_924 ();
 FILLCELL_X1 FILLER_0_72_942 ();
 FILLCELL_X1 FILLER_0_72_953 ();
 FILLCELL_X1 FILLER_0_72_979 ();
 FILLCELL_X2 FILLER_0_72_1053 ();
 FILLCELL_X4 FILLER_0_72_1059 ();
 FILLCELL_X1 FILLER_0_72_1063 ();
 FILLCELL_X8 FILLER_0_72_1067 ();
 FILLCELL_X1 FILLER_0_72_1075 ();
 FILLCELL_X2 FILLER_0_72_1084 ();
 FILLCELL_X1 FILLER_0_72_1086 ();
 FILLCELL_X2 FILLER_0_72_1094 ();
 FILLCELL_X1 FILLER_0_72_1096 ();
 FILLCELL_X32 FILLER_0_73_1 ();
 FILLCELL_X32 FILLER_0_73_33 ();
 FILLCELL_X32 FILLER_0_73_65 ();
 FILLCELL_X32 FILLER_0_73_97 ();
 FILLCELL_X32 FILLER_0_73_129 ();
 FILLCELL_X8 FILLER_0_73_161 ();
 FILLCELL_X4 FILLER_0_73_169 ();
 FILLCELL_X1 FILLER_0_73_173 ();
 FILLCELL_X1 FILLER_0_73_184 ();
 FILLCELL_X4 FILLER_0_73_194 ();
 FILLCELL_X2 FILLER_0_73_224 ();
 FILLCELL_X1 FILLER_0_73_226 ();
 FILLCELL_X4 FILLER_0_73_258 ();
 FILLCELL_X2 FILLER_0_73_335 ();
 FILLCELL_X1 FILLER_0_73_337 ();
 FILLCELL_X1 FILLER_0_73_378 ();
 FILLCELL_X8 FILLER_0_73_394 ();
 FILLCELL_X4 FILLER_0_73_402 ();
 FILLCELL_X8 FILLER_0_73_413 ();
 FILLCELL_X4 FILLER_0_73_421 ();
 FILLCELL_X1 FILLER_0_73_430 ();
 FILLCELL_X2 FILLER_0_73_438 ();
 FILLCELL_X1 FILLER_0_73_440 ();
 FILLCELL_X1 FILLER_0_73_451 ();
 FILLCELL_X4 FILLER_0_73_462 ();
 FILLCELL_X2 FILLER_0_73_466 ();
 FILLCELL_X2 FILLER_0_73_475 ();
 FILLCELL_X2 FILLER_0_73_549 ();
 FILLCELL_X2 FILLER_0_73_561 ();
 FILLCELL_X1 FILLER_0_73_563 ();
 FILLCELL_X1 FILLER_0_73_601 ();
 FILLCELL_X2 FILLER_0_73_612 ();
 FILLCELL_X1 FILLER_0_73_629 ();
 FILLCELL_X4 FILLER_0_73_647 ();
 FILLCELL_X2 FILLER_0_73_661 ();
 FILLCELL_X1 FILLER_0_73_663 ();
 FILLCELL_X2 FILLER_0_73_699 ();
 FILLCELL_X1 FILLER_0_73_701 ();
 FILLCELL_X1 FILLER_0_73_719 ();
 FILLCELL_X2 FILLER_0_73_747 ();
 FILLCELL_X2 FILLER_0_73_759 ();
 FILLCELL_X2 FILLER_0_73_796 ();
 FILLCELL_X1 FILLER_0_73_823 ();
 FILLCELL_X2 FILLER_0_73_834 ();
 FILLCELL_X4 FILLER_0_73_843 ();
 FILLCELL_X1 FILLER_0_73_847 ();
 FILLCELL_X2 FILLER_0_73_880 ();
 FILLCELL_X2 FILLER_0_73_902 ();
 FILLCELL_X1 FILLER_0_73_919 ();
 FILLCELL_X2 FILLER_0_73_957 ();
 FILLCELL_X1 FILLER_0_73_959 ();
 FILLCELL_X2 FILLER_0_73_980 ();
 FILLCELL_X4 FILLER_0_73_1050 ();
 FILLCELL_X2 FILLER_0_73_1054 ();
 FILLCELL_X1 FILLER_0_73_1056 ();
 FILLCELL_X2 FILLER_0_73_1106 ();
 FILLCELL_X2 FILLER_0_73_1124 ();
 FILLCELL_X2 FILLER_0_73_1146 ();
 FILLCELL_X32 FILLER_0_74_1 ();
 FILLCELL_X32 FILLER_0_74_33 ();
 FILLCELL_X32 FILLER_0_74_65 ();
 FILLCELL_X32 FILLER_0_74_97 ();
 FILLCELL_X32 FILLER_0_74_129 ();
 FILLCELL_X8 FILLER_0_74_161 ();
 FILLCELL_X1 FILLER_0_74_169 ();
 FILLCELL_X4 FILLER_0_74_185 ();
 FILLCELL_X2 FILLER_0_74_244 ();
 FILLCELL_X1 FILLER_0_74_246 ();
 FILLCELL_X1 FILLER_0_74_254 ();
 FILLCELL_X2 FILLER_0_74_289 ();
 FILLCELL_X4 FILLER_0_74_328 ();
 FILLCELL_X2 FILLER_0_74_365 ();
 FILLCELL_X4 FILLER_0_74_377 ();
 FILLCELL_X1 FILLER_0_74_381 ();
 FILLCELL_X4 FILLER_0_74_388 ();
 FILLCELL_X1 FILLER_0_74_392 ();
 FILLCELL_X2 FILLER_0_74_403 ();
 FILLCELL_X1 FILLER_0_74_405 ();
 FILLCELL_X2 FILLER_0_74_441 ();
 FILLCELL_X1 FILLER_0_74_443 ();
 FILLCELL_X2 FILLER_0_74_463 ();
 FILLCELL_X8 FILLER_0_74_476 ();
 FILLCELL_X1 FILLER_0_74_484 ();
 FILLCELL_X1 FILLER_0_74_575 ();
 FILLCELL_X2 FILLER_0_74_618 ();
 FILLCELL_X1 FILLER_0_74_620 ();
 FILLCELL_X1 FILLER_0_74_656 ();
 FILLCELL_X4 FILLER_0_74_674 ();
 FILLCELL_X2 FILLER_0_74_715 ();
 FILLCELL_X1 FILLER_0_74_724 ();
 FILLCELL_X1 FILLER_0_74_735 ();
 FILLCELL_X2 FILLER_0_74_760 ();
 FILLCELL_X1 FILLER_0_74_797 ();
 FILLCELL_X2 FILLER_0_74_815 ();
 FILLCELL_X1 FILLER_0_74_817 ();
 FILLCELL_X8 FILLER_0_74_833 ();
 FILLCELL_X1 FILLER_0_74_873 ();
 FILLCELL_X2 FILLER_0_74_908 ();
 FILLCELL_X1 FILLER_0_74_946 ();
 FILLCELL_X2 FILLER_0_74_990 ();
 FILLCELL_X1 FILLER_0_74_1007 ();
 FILLCELL_X8 FILLER_0_74_1042 ();
 FILLCELL_X2 FILLER_0_74_1050 ();
 FILLCELL_X1 FILLER_0_74_1052 ();
 FILLCELL_X2 FILLER_0_74_1126 ();
 FILLCELL_X8 FILLER_0_74_1135 ();
 FILLCELL_X4 FILLER_0_74_1143 ();
 FILLCELL_X1 FILLER_0_74_1147 ();
 FILLCELL_X16 FILLER_0_75_1 ();
 FILLCELL_X8 FILLER_0_75_17 ();
 FILLCELL_X4 FILLER_0_75_25 ();
 FILLCELL_X2 FILLER_0_75_29 ();
 FILLCELL_X1 FILLER_0_75_31 ();
 FILLCELL_X32 FILLER_0_75_57 ();
 FILLCELL_X32 FILLER_0_75_89 ();
 FILLCELL_X32 FILLER_0_75_121 ();
 FILLCELL_X16 FILLER_0_75_153 ();
 FILLCELL_X4 FILLER_0_75_169 ();
 FILLCELL_X2 FILLER_0_75_173 ();
 FILLCELL_X1 FILLER_0_75_175 ();
 FILLCELL_X4 FILLER_0_75_196 ();
 FILLCELL_X1 FILLER_0_75_205 ();
 FILLCELL_X1 FILLER_0_75_260 ();
 FILLCELL_X1 FILLER_0_75_293 ();
 FILLCELL_X1 FILLER_0_75_323 ();
 FILLCELL_X1 FILLER_0_75_374 ();
 FILLCELL_X4 FILLER_0_75_385 ();
 FILLCELL_X2 FILLER_0_75_396 ();
 FILLCELL_X1 FILLER_0_75_398 ();
 FILLCELL_X2 FILLER_0_75_409 ();
 FILLCELL_X1 FILLER_0_75_411 ();
 FILLCELL_X1 FILLER_0_75_417 ();
 FILLCELL_X4 FILLER_0_75_430 ();
 FILLCELL_X2 FILLER_0_75_444 ();
 FILLCELL_X8 FILLER_0_75_460 ();
 FILLCELL_X2 FILLER_0_75_468 ();
 FILLCELL_X4 FILLER_0_75_480 ();
 FILLCELL_X1 FILLER_0_75_484 ();
 FILLCELL_X2 FILLER_0_75_492 ();
 FILLCELL_X2 FILLER_0_75_504 ();
 FILLCELL_X4 FILLER_0_75_526 ();
 FILLCELL_X1 FILLER_0_75_549 ();
 FILLCELL_X2 FILLER_0_75_651 ();
 FILLCELL_X1 FILLER_0_75_668 ();
 FILLCELL_X2 FILLER_0_75_696 ();
 FILLCELL_X1 FILLER_0_75_738 ();
 FILLCELL_X1 FILLER_0_75_759 ();
 FILLCELL_X2 FILLER_0_75_774 ();
 FILLCELL_X1 FILLER_0_75_841 ();
 FILLCELL_X2 FILLER_0_75_847 ();
 FILLCELL_X1 FILLER_0_75_849 ();
 FILLCELL_X2 FILLER_0_75_860 ();
 FILLCELL_X1 FILLER_0_75_879 ();
 FILLCELL_X1 FILLER_0_75_897 ();
 FILLCELL_X2 FILLER_0_75_932 ();
 FILLCELL_X1 FILLER_0_75_966 ();
 FILLCELL_X1 FILLER_0_75_977 ();
 FILLCELL_X1 FILLER_0_75_1003 ();
 FILLCELL_X2 FILLER_0_75_1014 ();
 FILLCELL_X1 FILLER_0_75_1016 ();
 FILLCELL_X4 FILLER_0_75_1031 ();
 FILLCELL_X2 FILLER_0_75_1035 ();
 FILLCELL_X1 FILLER_0_75_1037 ();
 FILLCELL_X1 FILLER_0_75_1061 ();
 FILLCELL_X2 FILLER_0_75_1073 ();
 FILLCELL_X1 FILLER_0_75_1095 ();
 FILLCELL_X1 FILLER_0_75_1147 ();
 FILLCELL_X32 FILLER_0_76_1 ();
 FILLCELL_X32 FILLER_0_76_33 ();
 FILLCELL_X32 FILLER_0_76_65 ();
 FILLCELL_X32 FILLER_0_76_97 ();
 FILLCELL_X32 FILLER_0_76_129 ();
 FILLCELL_X4 FILLER_0_76_161 ();
 FILLCELL_X2 FILLER_0_76_165 ();
 FILLCELL_X4 FILLER_0_76_228 ();
 FILLCELL_X2 FILLER_0_76_232 ();
 FILLCELL_X1 FILLER_0_76_265 ();
 FILLCELL_X1 FILLER_0_76_283 ();
 FILLCELL_X2 FILLER_0_76_333 ();
 FILLCELL_X1 FILLER_0_76_335 ();
 FILLCELL_X2 FILLER_0_76_346 ();
 FILLCELL_X1 FILLER_0_76_348 ();
 FILLCELL_X2 FILLER_0_76_411 ();
 FILLCELL_X4 FILLER_0_76_423 ();
 FILLCELL_X1 FILLER_0_76_427 ();
 FILLCELL_X2 FILLER_0_76_440 ();
 FILLCELL_X4 FILLER_0_76_469 ();
 FILLCELL_X2 FILLER_0_76_490 ();
 FILLCELL_X1 FILLER_0_76_492 ();
 FILLCELL_X1 FILLER_0_76_503 ();
 FILLCELL_X1 FILLER_0_76_514 ();
 FILLCELL_X4 FILLER_0_76_535 ();
 FILLCELL_X2 FILLER_0_76_557 ();
 FILLCELL_X2 FILLER_0_76_591 ();
 FILLCELL_X1 FILLER_0_76_613 ();
 FILLCELL_X2 FILLER_0_76_645 ();
 FILLCELL_X1 FILLER_0_76_647 ();
 FILLCELL_X1 FILLER_0_76_701 ();
 FILLCELL_X8 FILLER_0_76_752 ();
 FILLCELL_X2 FILLER_0_76_760 ();
 FILLCELL_X8 FILLER_0_76_793 ();
 FILLCELL_X1 FILLER_0_76_801 ();
 FILLCELL_X4 FILLER_0_76_807 ();
 FILLCELL_X1 FILLER_0_76_811 ();
 FILLCELL_X2 FILLER_0_76_827 ();
 FILLCELL_X2 FILLER_0_76_874 ();
 FILLCELL_X1 FILLER_0_76_876 ();
 FILLCELL_X2 FILLER_0_76_894 ();
 FILLCELL_X1 FILLER_0_76_896 ();
 FILLCELL_X2 FILLER_0_76_917 ();
 FILLCELL_X2 FILLER_0_76_960 ();
 FILLCELL_X1 FILLER_0_76_962 ();
 FILLCELL_X2 FILLER_0_76_980 ();
 FILLCELL_X1 FILLER_0_76_982 ();
 FILLCELL_X2 FILLER_0_76_1023 ();
 FILLCELL_X4 FILLER_0_76_1035 ();
 FILLCELL_X2 FILLER_0_76_1039 ();
 FILLCELL_X1 FILLER_0_76_1041 ();
 FILLCELL_X1 FILLER_0_76_1094 ();
 FILLCELL_X2 FILLER_0_76_1132 ();
 FILLCELL_X32 FILLER_0_77_1 ();
 FILLCELL_X32 FILLER_0_77_33 ();
 FILLCELL_X32 FILLER_0_77_65 ();
 FILLCELL_X32 FILLER_0_77_97 ();
 FILLCELL_X32 FILLER_0_77_129 ();
 FILLCELL_X8 FILLER_0_77_161 ();
 FILLCELL_X4 FILLER_0_77_169 ();
 FILLCELL_X2 FILLER_0_77_173 ();
 FILLCELL_X1 FILLER_0_77_175 ();
 FILLCELL_X4 FILLER_0_77_186 ();
 FILLCELL_X2 FILLER_0_77_190 ();
 FILLCELL_X1 FILLER_0_77_259 ();
 FILLCELL_X1 FILLER_0_77_270 ();
 FILLCELL_X2 FILLER_0_77_313 ();
 FILLCELL_X1 FILLER_0_77_315 ();
 FILLCELL_X1 FILLER_0_77_377 ();
 FILLCELL_X2 FILLER_0_77_388 ();
 FILLCELL_X1 FILLER_0_77_390 ();
 FILLCELL_X1 FILLER_0_77_393 ();
 FILLCELL_X8 FILLER_0_77_407 ();
 FILLCELL_X2 FILLER_0_77_415 ();
 FILLCELL_X8 FILLER_0_77_427 ();
 FILLCELL_X4 FILLER_0_77_435 ();
 FILLCELL_X2 FILLER_0_77_439 ();
 FILLCELL_X2 FILLER_0_77_466 ();
 FILLCELL_X2 FILLER_0_77_479 ();
 FILLCELL_X1 FILLER_0_77_481 ();
 FILLCELL_X1 FILLER_0_77_503 ();
 FILLCELL_X1 FILLER_0_77_509 ();
 FILLCELL_X1 FILLER_0_77_520 ();
 FILLCELL_X2 FILLER_0_77_541 ();
 FILLCELL_X1 FILLER_0_77_543 ();
 FILLCELL_X2 FILLER_0_77_561 ();
 FILLCELL_X1 FILLER_0_77_563 ();
 FILLCELL_X1 FILLER_0_77_569 ();
 FILLCELL_X1 FILLER_0_77_580 ();
 FILLCELL_X1 FILLER_0_77_596 ();
 FILLCELL_X1 FILLER_0_77_612 ();
 FILLCELL_X1 FILLER_0_77_637 ();
 FILLCELL_X2 FILLER_0_77_662 ();
 FILLCELL_X1 FILLER_0_77_709 ();
 FILLCELL_X2 FILLER_0_77_720 ();
 FILLCELL_X1 FILLER_0_77_732 ();
 FILLCELL_X4 FILLER_0_77_747 ();
 FILLCELL_X2 FILLER_0_77_751 ();
 FILLCELL_X1 FILLER_0_77_753 ();
 FILLCELL_X4 FILLER_0_77_793 ();
 FILLCELL_X2 FILLER_0_77_797 ();
 FILLCELL_X2 FILLER_0_77_809 ();
 FILLCELL_X2 FILLER_0_77_816 ();
 FILLCELL_X1 FILLER_0_77_818 ();
 FILLCELL_X1 FILLER_0_77_829 ();
 FILLCELL_X2 FILLER_0_77_840 ();
 FILLCELL_X1 FILLER_0_77_842 ();
 FILLCELL_X1 FILLER_0_77_868 ();
 FILLCELL_X2 FILLER_0_77_886 ();
 FILLCELL_X1 FILLER_0_77_888 ();
 FILLCELL_X2 FILLER_0_77_906 ();
 FILLCELL_X2 FILLER_0_77_940 ();
 FILLCELL_X1 FILLER_0_77_942 ();
 FILLCELL_X2 FILLER_0_77_960 ();
 FILLCELL_X2 FILLER_0_77_972 ();
 FILLCELL_X1 FILLER_0_77_991 ();
 FILLCELL_X1 FILLER_0_77_1012 ();
 FILLCELL_X2 FILLER_0_77_1028 ();
 FILLCELL_X1 FILLER_0_77_1030 ();
 FILLCELL_X2 FILLER_0_77_1046 ();
 FILLCELL_X1 FILLER_0_77_1048 ();
 FILLCELL_X8 FILLER_0_77_1072 ();
 FILLCELL_X1 FILLER_0_77_1080 ();
 FILLCELL_X2 FILLER_0_77_1146 ();
 FILLCELL_X32 FILLER_0_78_1 ();
 FILLCELL_X32 FILLER_0_78_33 ();
 FILLCELL_X32 FILLER_0_78_65 ();
 FILLCELL_X32 FILLER_0_78_97 ();
 FILLCELL_X32 FILLER_0_78_129 ();
 FILLCELL_X8 FILLER_0_78_161 ();
 FILLCELL_X4 FILLER_0_78_198 ();
 FILLCELL_X4 FILLER_0_78_212 ();
 FILLCELL_X4 FILLER_0_78_226 ();
 FILLCELL_X4 FILLER_0_78_240 ();
 FILLCELL_X1 FILLER_0_78_262 ();
 FILLCELL_X1 FILLER_0_78_277 ();
 FILLCELL_X2 FILLER_0_78_295 ();
 FILLCELL_X2 FILLER_0_78_306 ();
 FILLCELL_X1 FILLER_0_78_317 ();
 FILLCELL_X2 FILLER_0_78_342 ();
 FILLCELL_X2 FILLER_0_78_354 ();
 FILLCELL_X1 FILLER_0_78_356 ();
 FILLCELL_X2 FILLER_0_78_401 ();
 FILLCELL_X1 FILLER_0_78_417 ();
 FILLCELL_X2 FILLER_0_78_439 ();
 FILLCELL_X1 FILLER_0_78_441 ();
 FILLCELL_X8 FILLER_0_78_456 ();
 FILLCELL_X4 FILLER_0_78_464 ();
 FILLCELL_X1 FILLER_0_78_513 ();
 FILLCELL_X2 FILLER_0_78_524 ();
 FILLCELL_X2 FILLER_0_78_569 ();
 FILLCELL_X1 FILLER_0_78_571 ();
 FILLCELL_X2 FILLER_0_78_596 ();
 FILLCELL_X1 FILLER_0_78_598 ();
 FILLCELL_X2 FILLER_0_78_606 ();
 FILLCELL_X2 FILLER_0_78_629 ();
 FILLCELL_X1 FILLER_0_78_632 ();
 FILLCELL_X2 FILLER_0_78_675 ();
 FILLCELL_X1 FILLER_0_78_677 ();
 FILLCELL_X1 FILLER_0_78_688 ();
 FILLCELL_X2 FILLER_0_78_706 ();
 FILLCELL_X1 FILLER_0_78_708 ();
 FILLCELL_X2 FILLER_0_78_731 ();
 FILLCELL_X1 FILLER_0_78_743 ();
 FILLCELL_X4 FILLER_0_78_758 ();
 FILLCELL_X1 FILLER_0_78_762 ();
 FILLCELL_X8 FILLER_0_78_770 ();
 FILLCELL_X2 FILLER_0_78_778 ();
 FILLCELL_X1 FILLER_0_78_780 ();
 FILLCELL_X8 FILLER_0_78_785 ();
 FILLCELL_X4 FILLER_0_78_793 ();
 FILLCELL_X2 FILLER_0_78_797 ();
 FILLCELL_X1 FILLER_0_78_799 ();
 FILLCELL_X4 FILLER_0_78_810 ();
 FILLCELL_X1 FILLER_0_78_846 ();
 FILLCELL_X4 FILLER_0_78_906 ();
 FILLCELL_X2 FILLER_0_78_932 ();
 FILLCELL_X2 FILLER_0_78_961 ();
 FILLCELL_X1 FILLER_0_78_963 ();
 FILLCELL_X2 FILLER_0_78_981 ();
 FILLCELL_X1 FILLER_0_78_983 ();
 FILLCELL_X2 FILLER_0_78_994 ();
 FILLCELL_X1 FILLER_0_78_996 ();
 FILLCELL_X4 FILLER_0_78_1019 ();
 FILLCELL_X16 FILLER_0_78_1033 ();
 FILLCELL_X8 FILLER_0_78_1049 ();
 FILLCELL_X1 FILLER_0_78_1057 ();
 FILLCELL_X2 FILLER_0_78_1068 ();
 FILLCELL_X2 FILLER_0_78_1073 ();
 FILLCELL_X4 FILLER_0_78_1098 ();
 FILLCELL_X1 FILLER_0_78_1105 ();
 FILLCELL_X4 FILLER_0_78_1143 ();
 FILLCELL_X1 FILLER_0_78_1147 ();
 FILLCELL_X32 FILLER_0_79_1 ();
 FILLCELL_X32 FILLER_0_79_33 ();
 FILLCELL_X32 FILLER_0_79_65 ();
 FILLCELL_X32 FILLER_0_79_97 ();
 FILLCELL_X16 FILLER_0_79_129 ();
 FILLCELL_X8 FILLER_0_79_145 ();
 FILLCELL_X4 FILLER_0_79_153 ();
 FILLCELL_X2 FILLER_0_79_157 ();
 FILLCELL_X4 FILLER_0_79_174 ();
 FILLCELL_X1 FILLER_0_79_178 ();
 FILLCELL_X2 FILLER_0_79_189 ();
 FILLCELL_X4 FILLER_0_79_218 ();
 FILLCELL_X4 FILLER_0_79_273 ();
 FILLCELL_X1 FILLER_0_79_291 ();
 FILLCELL_X2 FILLER_0_79_317 ();
 FILLCELL_X1 FILLER_0_79_319 ();
 FILLCELL_X2 FILLER_0_79_347 ();
 FILLCELL_X1 FILLER_0_79_378 ();
 FILLCELL_X2 FILLER_0_79_404 ();
 FILLCELL_X8 FILLER_0_79_413 ();
 FILLCELL_X1 FILLER_0_79_421 ();
 FILLCELL_X4 FILLER_0_79_434 ();
 FILLCELL_X2 FILLER_0_79_438 ();
 FILLCELL_X4 FILLER_0_79_450 ();
 FILLCELL_X1 FILLER_0_79_454 ();
 FILLCELL_X8 FILLER_0_79_471 ();
 FILLCELL_X4 FILLER_0_79_479 ();
 FILLCELL_X8 FILLER_0_79_516 ();
 FILLCELL_X1 FILLER_0_79_585 ();
 FILLCELL_X1 FILLER_0_79_596 ();
 FILLCELL_X2 FILLER_0_79_607 ();
 FILLCELL_X1 FILLER_0_79_609 ();
 FILLCELL_X2 FILLER_0_79_623 ();
 FILLCELL_X1 FILLER_0_79_696 ();
 FILLCELL_X1 FILLER_0_79_714 ();
 FILLCELL_X8 FILLER_0_79_792 ();
 FILLCELL_X4 FILLER_0_79_800 ();
 FILLCELL_X2 FILLER_0_79_804 ();
 FILLCELL_X2 FILLER_0_79_821 ();
 FILLCELL_X2 FILLER_0_79_854 ();
 FILLCELL_X1 FILLER_0_79_856 ();
 FILLCELL_X4 FILLER_0_79_867 ();
 FILLCELL_X1 FILLER_0_79_895 ();
 FILLCELL_X2 FILLER_0_79_906 ();
 FILLCELL_X1 FILLER_0_79_908 ();
 FILLCELL_X2 FILLER_0_79_933 ();
 FILLCELL_X1 FILLER_0_79_935 ();
 FILLCELL_X1 FILLER_0_79_951 ();
 FILLCELL_X1 FILLER_0_79_992 ();
 FILLCELL_X1 FILLER_0_79_1018 ();
 FILLCELL_X4 FILLER_0_79_1029 ();
 FILLCELL_X8 FILLER_0_79_1043 ();
 FILLCELL_X4 FILLER_0_79_1051 ();
 FILLCELL_X2 FILLER_0_79_1055 ();
 FILLCELL_X2 FILLER_0_79_1096 ();
 FILLCELL_X2 FILLER_0_79_1118 ();
 FILLCELL_X2 FILLER_0_79_1123 ();
 FILLCELL_X32 FILLER_0_80_1 ();
 FILLCELL_X32 FILLER_0_80_33 ();
 FILLCELL_X32 FILLER_0_80_65 ();
 FILLCELL_X32 FILLER_0_80_97 ();
 FILLCELL_X32 FILLER_0_80_129 ();
 FILLCELL_X2 FILLER_0_80_161 ();
 FILLCELL_X1 FILLER_0_80_173 ();
 FILLCELL_X1 FILLER_0_80_183 ();
 FILLCELL_X1 FILLER_0_80_189 ();
 FILLCELL_X2 FILLER_0_80_200 ();
 FILLCELL_X1 FILLER_0_80_202 ();
 FILLCELL_X1 FILLER_0_80_225 ();
 FILLCELL_X1 FILLER_0_80_261 ();
 FILLCELL_X1 FILLER_0_80_286 ();
 FILLCELL_X1 FILLER_0_80_299 ();
 FILLCELL_X2 FILLER_0_80_331 ();
 FILLCELL_X2 FILLER_0_80_340 ();
 FILLCELL_X1 FILLER_0_80_352 ();
 FILLCELL_X1 FILLER_0_80_368 ();
 FILLCELL_X1 FILLER_0_80_379 ();
 FILLCELL_X1 FILLER_0_80_395 ();
 FILLCELL_X1 FILLER_0_80_413 ();
 FILLCELL_X16 FILLER_0_80_442 ();
 FILLCELL_X1 FILLER_0_80_458 ();
 FILLCELL_X1 FILLER_0_80_461 ();
 FILLCELL_X8 FILLER_0_80_472 ();
 FILLCELL_X4 FILLER_0_80_480 ();
 FILLCELL_X2 FILLER_0_80_502 ();
 FILLCELL_X1 FILLER_0_80_504 ();
 FILLCELL_X1 FILLER_0_80_522 ();
 FILLCELL_X1 FILLER_0_80_533 ();
 FILLCELL_X4 FILLER_0_80_551 ();
 FILLCELL_X1 FILLER_0_80_575 ();
 FILLCELL_X4 FILLER_0_80_608 ();
 FILLCELL_X1 FILLER_0_80_612 ();
 FILLCELL_X2 FILLER_0_80_628 ();
 FILLCELL_X1 FILLER_0_80_630 ();
 FILLCELL_X1 FILLER_0_80_632 ();
 FILLCELL_X2 FILLER_0_80_668 ();
 FILLCELL_X2 FILLER_0_80_741 ();
 FILLCELL_X16 FILLER_0_80_748 ();
 FILLCELL_X4 FILLER_0_80_764 ();
 FILLCELL_X1 FILLER_0_80_768 ();
 FILLCELL_X1 FILLER_0_80_772 ();
 FILLCELL_X8 FILLER_0_80_783 ();
 FILLCELL_X16 FILLER_0_80_801 ();
 FILLCELL_X2 FILLER_0_80_817 ();
 FILLCELL_X1 FILLER_0_80_819 ();
 FILLCELL_X2 FILLER_0_80_840 ();
 FILLCELL_X2 FILLER_0_80_861 ();
 FILLCELL_X1 FILLER_0_80_863 ();
 FILLCELL_X4 FILLER_0_80_932 ();
 FILLCELL_X4 FILLER_0_80_961 ();
 FILLCELL_X2 FILLER_0_80_975 ();
 FILLCELL_X1 FILLER_0_80_977 ();
 FILLCELL_X8 FILLER_0_80_1030 ();
 FILLCELL_X2 FILLER_0_80_1038 ();
 FILLCELL_X1 FILLER_0_80_1080 ();
 FILLCELL_X2 FILLER_0_80_1089 ();
 FILLCELL_X1 FILLER_0_80_1091 ();
 FILLCELL_X2 FILLER_0_80_1096 ();
 FILLCELL_X1 FILLER_0_80_1098 ();
 FILLCELL_X1 FILLER_0_80_1103 ();
 FILLCELL_X1 FILLER_0_80_1147 ();
 FILLCELL_X32 FILLER_0_81_1 ();
 FILLCELL_X32 FILLER_0_81_33 ();
 FILLCELL_X32 FILLER_0_81_65 ();
 FILLCELL_X32 FILLER_0_81_97 ();
 FILLCELL_X32 FILLER_0_81_129 ();
 FILLCELL_X16 FILLER_0_81_161 ();
 FILLCELL_X8 FILLER_0_81_177 ();
 FILLCELL_X1 FILLER_0_81_185 ();
 FILLCELL_X1 FILLER_0_81_201 ();
 FILLCELL_X2 FILLER_0_81_234 ();
 FILLCELL_X1 FILLER_0_81_236 ();
 FILLCELL_X1 FILLER_0_81_273 ();
 FILLCELL_X1 FILLER_0_81_289 ();
 FILLCELL_X1 FILLER_0_81_310 ();
 FILLCELL_X2 FILLER_0_81_453 ();
 FILLCELL_X8 FILLER_0_81_458 ();
 FILLCELL_X1 FILLER_0_81_469 ();
 FILLCELL_X2 FILLER_0_81_522 ();
 FILLCELL_X4 FILLER_0_81_540 ();
 FILLCELL_X2 FILLER_0_81_549 ();
 FILLCELL_X1 FILLER_0_81_574 ();
 FILLCELL_X2 FILLER_0_81_602 ();
 FILLCELL_X1 FILLER_0_81_604 ();
 FILLCELL_X1 FILLER_0_81_617 ();
 FILLCELL_X2 FILLER_0_81_653 ();
 FILLCELL_X1 FILLER_0_81_655 ();
 FILLCELL_X1 FILLER_0_81_679 ();
 FILLCELL_X1 FILLER_0_81_723 ();
 FILLCELL_X16 FILLER_0_81_741 ();
 FILLCELL_X1 FILLER_0_81_764 ();
 FILLCELL_X4 FILLER_0_81_769 ();
 FILLCELL_X2 FILLER_0_81_780 ();
 FILLCELL_X2 FILLER_0_81_788 ();
 FILLCELL_X2 FILLER_0_81_800 ();
 FILLCELL_X1 FILLER_0_81_817 ();
 FILLCELL_X1 FILLER_0_81_822 ();
 FILLCELL_X1 FILLER_0_81_828 ();
 FILLCELL_X2 FILLER_0_81_849 ();
 FILLCELL_X1 FILLER_0_81_883 ();
 FILLCELL_X2 FILLER_0_81_894 ();
 FILLCELL_X1 FILLER_0_81_896 ();
 FILLCELL_X2 FILLER_0_81_924 ();
 FILLCELL_X4 FILLER_0_81_1021 ();
 FILLCELL_X1 FILLER_0_81_1065 ();
 FILLCELL_X1 FILLER_0_81_1070 ();
 FILLCELL_X1 FILLER_0_81_1075 ();
 FILLCELL_X1 FILLER_0_81_1084 ();
 FILLCELL_X1 FILLER_0_81_1087 ();
 FILLCELL_X1 FILLER_0_81_1112 ();
 FILLCELL_X2 FILLER_0_81_1117 ();
 FILLCELL_X2 FILLER_0_81_1123 ();
 FILLCELL_X1 FILLER_0_81_1125 ();
 FILLCELL_X2 FILLER_0_81_1146 ();
 FILLCELL_X32 FILLER_0_82_1 ();
 FILLCELL_X32 FILLER_0_82_33 ();
 FILLCELL_X32 FILLER_0_82_65 ();
 FILLCELL_X32 FILLER_0_82_97 ();
 FILLCELL_X32 FILLER_0_82_129 ();
 FILLCELL_X16 FILLER_0_82_161 ();
 FILLCELL_X4 FILLER_0_82_177 ();
 FILLCELL_X2 FILLER_0_82_181 ();
 FILLCELL_X4 FILLER_0_82_198 ();
 FILLCELL_X2 FILLER_0_82_207 ();
 FILLCELL_X1 FILLER_0_82_209 ();
 FILLCELL_X1 FILLER_0_82_223 ();
 FILLCELL_X8 FILLER_0_82_230 ();
 FILLCELL_X2 FILLER_0_82_238 ();
 FILLCELL_X1 FILLER_0_82_240 ();
 FILLCELL_X2 FILLER_0_82_255 ();
 FILLCELL_X4 FILLER_0_82_267 ();
 FILLCELL_X16 FILLER_0_82_368 ();
 FILLCELL_X8 FILLER_0_82_384 ();
 FILLCELL_X8 FILLER_0_82_471 ();
 FILLCELL_X4 FILLER_0_82_479 ();
 FILLCELL_X8 FILLER_0_82_486 ();
 FILLCELL_X1 FILLER_0_82_494 ();
 FILLCELL_X1 FILLER_0_82_498 ();
 FILLCELL_X4 FILLER_0_82_540 ();
 FILLCELL_X4 FILLER_0_82_551 ();
 FILLCELL_X2 FILLER_0_82_555 ();
 FILLCELL_X1 FILLER_0_82_557 ();
 FILLCELL_X2 FILLER_0_82_568 ();
 FILLCELL_X1 FILLER_0_82_575 ();
 FILLCELL_X2 FILLER_0_82_591 ();
 FILLCELL_X1 FILLER_0_82_593 ();
 FILLCELL_X2 FILLER_0_82_624 ();
 FILLCELL_X2 FILLER_0_82_642 ();
 FILLCELL_X2 FILLER_0_82_654 ();
 FILLCELL_X2 FILLER_0_82_661 ();
 FILLCELL_X1 FILLER_0_82_695 ();
 FILLCELL_X2 FILLER_0_82_709 ();
 FILLCELL_X1 FILLER_0_82_711 ();
 FILLCELL_X1 FILLER_0_82_723 ();
 FILLCELL_X2 FILLER_0_82_752 ();
 FILLCELL_X1 FILLER_0_82_754 ();
 FILLCELL_X2 FILLER_0_82_779 ();
 FILLCELL_X1 FILLER_0_82_781 ();
 FILLCELL_X2 FILLER_0_82_792 ();
 FILLCELL_X4 FILLER_0_82_804 ();
 FILLCELL_X2 FILLER_0_82_808 ();
 FILLCELL_X1 FILLER_0_82_829 ();
 FILLCELL_X4 FILLER_0_82_835 ();
 FILLCELL_X1 FILLER_0_82_839 ();
 FILLCELL_X4 FILLER_0_82_845 ();
 FILLCELL_X2 FILLER_0_82_849 ();
 FILLCELL_X4 FILLER_0_82_861 ();
 FILLCELL_X2 FILLER_0_82_865 ();
 FILLCELL_X1 FILLER_0_82_884 ();
 FILLCELL_X2 FILLER_0_82_902 ();
 FILLCELL_X1 FILLER_0_82_904 ();
 FILLCELL_X1 FILLER_0_82_920 ();
 FILLCELL_X1 FILLER_0_82_952 ();
 FILLCELL_X1 FILLER_0_82_963 ();
 FILLCELL_X2 FILLER_0_82_971 ();
 FILLCELL_X1 FILLER_0_82_973 ();
 FILLCELL_X4 FILLER_0_82_1004 ();
 FILLCELL_X8 FILLER_0_82_1028 ();
 FILLCELL_X2 FILLER_0_82_1036 ();
 FILLCELL_X8 FILLER_0_82_1041 ();
 FILLCELL_X4 FILLER_0_82_1049 ();
 FILLCELL_X1 FILLER_0_82_1053 ();
 FILLCELL_X1 FILLER_0_82_1070 ();
 FILLCELL_X1 FILLER_0_82_1125 ();
 FILLCELL_X2 FILLER_0_82_1146 ();
 FILLCELL_X32 FILLER_0_83_1 ();
 FILLCELL_X32 FILLER_0_83_33 ();
 FILLCELL_X32 FILLER_0_83_65 ();
 FILLCELL_X32 FILLER_0_83_97 ();
 FILLCELL_X32 FILLER_0_83_129 ();
 FILLCELL_X8 FILLER_0_83_161 ();
 FILLCELL_X4 FILLER_0_83_169 ();
 FILLCELL_X4 FILLER_0_83_238 ();
 FILLCELL_X1 FILLER_0_83_297 ();
 FILLCELL_X2 FILLER_0_83_364 ();
 FILLCELL_X1 FILLER_0_83_370 ();
 FILLCELL_X2 FILLER_0_83_378 ();
 FILLCELL_X2 FILLER_0_83_390 ();
 FILLCELL_X2 FILLER_0_83_395 ();
 FILLCELL_X1 FILLER_0_83_408 ();
 FILLCELL_X1 FILLER_0_83_455 ();
 FILLCELL_X8 FILLER_0_83_475 ();
 FILLCELL_X1 FILLER_0_83_483 ();
 FILLCELL_X1 FILLER_0_83_498 ();
 FILLCELL_X8 FILLER_0_83_522 ();
 FILLCELL_X2 FILLER_0_83_565 ();
 FILLCELL_X1 FILLER_0_83_567 ();
 FILLCELL_X4 FILLER_0_83_588 ();
 FILLCELL_X2 FILLER_0_83_592 ();
 FILLCELL_X4 FILLER_0_83_644 ();
 FILLCELL_X2 FILLER_0_83_648 ();
 FILLCELL_X1 FILLER_0_83_650 ();
 FILLCELL_X1 FILLER_0_83_671 ();
 FILLCELL_X2 FILLER_0_83_704 ();
 FILLCELL_X2 FILLER_0_83_740 ();
 FILLCELL_X2 FILLER_0_83_752 ();
 FILLCELL_X2 FILLER_0_83_764 ();
 FILLCELL_X2 FILLER_0_83_790 ();
 FILLCELL_X16 FILLER_0_83_795 ();
 FILLCELL_X4 FILLER_0_83_811 ();
 FILLCELL_X1 FILLER_0_83_815 ();
 FILLCELL_X1 FILLER_0_83_841 ();
 FILLCELL_X1 FILLER_0_83_852 ();
 FILLCELL_X1 FILLER_0_83_858 ();
 FILLCELL_X1 FILLER_0_83_869 ();
 FILLCELL_X4 FILLER_0_83_887 ();
 FILLCELL_X1 FILLER_0_83_901 ();
 FILLCELL_X2 FILLER_0_83_912 ();
 FILLCELL_X2 FILLER_0_83_924 ();
 FILLCELL_X2 FILLER_0_83_936 ();
 FILLCELL_X1 FILLER_0_83_952 ();
 FILLCELL_X2 FILLER_0_83_977 ();
 FILLCELL_X4 FILLER_0_83_989 ();
 FILLCELL_X2 FILLER_0_83_1002 ();
 FILLCELL_X1 FILLER_0_83_1004 ();
 FILLCELL_X2 FILLER_0_83_1014 ();
 FILLCELL_X1 FILLER_0_83_1016 ();
 FILLCELL_X32 FILLER_0_83_1022 ();
 FILLCELL_X2 FILLER_0_83_1054 ();
 FILLCELL_X2 FILLER_0_83_1100 ();
 FILLCELL_X1 FILLER_0_83_1112 ();
 FILLCELL_X1 FILLER_0_83_1120 ();
 FILLCELL_X2 FILLER_0_83_1132 ();
 FILLCELL_X32 FILLER_0_84_1 ();
 FILLCELL_X32 FILLER_0_84_33 ();
 FILLCELL_X32 FILLER_0_84_65 ();
 FILLCELL_X32 FILLER_0_84_97 ();
 FILLCELL_X32 FILLER_0_84_129 ();
 FILLCELL_X16 FILLER_0_84_161 ();
 FILLCELL_X4 FILLER_0_84_177 ();
 FILLCELL_X2 FILLER_0_84_181 ();
 FILLCELL_X1 FILLER_0_84_183 ();
 FILLCELL_X8 FILLER_0_84_194 ();
 FILLCELL_X2 FILLER_0_84_202 ();
 FILLCELL_X4 FILLER_0_84_219 ();
 FILLCELL_X1 FILLER_0_84_223 ();
 FILLCELL_X2 FILLER_0_84_254 ();
 FILLCELL_X1 FILLER_0_84_266 ();
 FILLCELL_X2 FILLER_0_84_272 ();
 FILLCELL_X1 FILLER_0_84_357 ();
 FILLCELL_X1 FILLER_0_84_371 ();
 FILLCELL_X1 FILLER_0_84_382 ();
 FILLCELL_X1 FILLER_0_84_390 ();
 FILLCELL_X2 FILLER_0_84_401 ();
 FILLCELL_X1 FILLER_0_84_403 ();
 FILLCELL_X2 FILLER_0_84_407 ();
 FILLCELL_X1 FILLER_0_84_409 ();
 FILLCELL_X1 FILLER_0_84_420 ();
 FILLCELL_X2 FILLER_0_84_448 ();
 FILLCELL_X2 FILLER_0_84_460 ();
 FILLCELL_X1 FILLER_0_84_462 ();
 FILLCELL_X4 FILLER_0_84_497 ();
 FILLCELL_X2 FILLER_0_84_501 ();
 FILLCELL_X8 FILLER_0_84_505 ();
 FILLCELL_X1 FILLER_0_84_516 ();
 FILLCELL_X2 FILLER_0_84_521 ();
 FILLCELL_X4 FILLER_0_84_574 ();
 FILLCELL_X16 FILLER_0_84_592 ();
 FILLCELL_X2 FILLER_0_84_608 ();
 FILLCELL_X2 FILLER_0_84_615 ();
 FILLCELL_X1 FILLER_0_84_617 ();
 FILLCELL_X2 FILLER_0_84_646 ();
 FILLCELL_X4 FILLER_0_84_683 ();
 FILLCELL_X1 FILLER_0_84_687 ();
 FILLCELL_X2 FILLER_0_84_761 ();
 FILLCELL_X4 FILLER_0_84_773 ();
 FILLCELL_X2 FILLER_0_84_777 ();
 FILLCELL_X1 FILLER_0_84_779 ();
 FILLCELL_X8 FILLER_0_84_811 ();
 FILLCELL_X4 FILLER_0_84_819 ();
 FILLCELL_X1 FILLER_0_84_823 ();
 FILLCELL_X4 FILLER_0_84_827 ();
 FILLCELL_X1 FILLER_0_84_871 ();
 FILLCELL_X2 FILLER_0_84_954 ();
 FILLCELL_X1 FILLER_0_84_956 ();
 FILLCELL_X2 FILLER_0_84_984 ();
 FILLCELL_X1 FILLER_0_84_986 ();
 FILLCELL_X2 FILLER_0_84_1011 ();
 FILLCELL_X4 FILLER_0_84_1028 ();
 FILLCELL_X1 FILLER_0_84_1073 ();
 FILLCELL_X1 FILLER_0_84_1105 ();
 FILLCELL_X8 FILLER_0_84_1126 ();
 FILLCELL_X4 FILLER_0_84_1134 ();
 FILLCELL_X2 FILLER_0_84_1145 ();
 FILLCELL_X1 FILLER_0_84_1147 ();
 FILLCELL_X32 FILLER_0_85_1 ();
 FILLCELL_X32 FILLER_0_85_33 ();
 FILLCELL_X32 FILLER_0_85_65 ();
 FILLCELL_X32 FILLER_0_85_97 ();
 FILLCELL_X32 FILLER_0_85_129 ();
 FILLCELL_X8 FILLER_0_85_161 ();
 FILLCELL_X4 FILLER_0_85_169 ();
 FILLCELL_X2 FILLER_0_85_212 ();
 FILLCELL_X2 FILLER_0_85_244 ();
 FILLCELL_X2 FILLER_0_85_286 ();
 FILLCELL_X4 FILLER_0_85_303 ();
 FILLCELL_X1 FILLER_0_85_307 ();
 FILLCELL_X1 FILLER_0_85_357 ();
 FILLCELL_X2 FILLER_0_85_371 ();
 FILLCELL_X1 FILLER_0_85_383 ();
 FILLCELL_X2 FILLER_0_85_394 ();
 FILLCELL_X1 FILLER_0_85_399 ();
 FILLCELL_X2 FILLER_0_85_414 ();
 FILLCELL_X2 FILLER_0_85_461 ();
 FILLCELL_X1 FILLER_0_85_463 ();
 FILLCELL_X2 FILLER_0_85_475 ();
 FILLCELL_X4 FILLER_0_85_494 ();
 FILLCELL_X2 FILLER_0_85_498 ();
 FILLCELL_X4 FILLER_0_85_534 ();
 FILLCELL_X2 FILLER_0_85_538 ();
 FILLCELL_X1 FILLER_0_85_540 ();
 FILLCELL_X2 FILLER_0_85_554 ();
 FILLCELL_X1 FILLER_0_85_569 ();
 FILLCELL_X1 FILLER_0_85_574 ();
 FILLCELL_X1 FILLER_0_85_579 ();
 FILLCELL_X1 FILLER_0_85_590 ();
 FILLCELL_X2 FILLER_0_85_596 ();
 FILLCELL_X1 FILLER_0_85_636 ();
 FILLCELL_X1 FILLER_0_85_642 ();
 FILLCELL_X2 FILLER_0_85_658 ();
 FILLCELL_X1 FILLER_0_85_660 ();
 FILLCELL_X4 FILLER_0_85_666 ();
 FILLCELL_X1 FILLER_0_85_670 ();
 FILLCELL_X4 FILLER_0_85_676 ();
 FILLCELL_X1 FILLER_0_85_680 ();
 FILLCELL_X2 FILLER_0_85_691 ();
 FILLCELL_X1 FILLER_0_85_693 ();
 FILLCELL_X4 FILLER_0_85_711 ();
 FILLCELL_X2 FILLER_0_85_715 ();
 FILLCELL_X2 FILLER_0_85_737 ();
 FILLCELL_X1 FILLER_0_85_739 ();
 FILLCELL_X8 FILLER_0_85_747 ();
 FILLCELL_X1 FILLER_0_85_755 ();
 FILLCELL_X4 FILLER_0_85_780 ();
 FILLCELL_X2 FILLER_0_85_784 ();
 FILLCELL_X1 FILLER_0_85_786 ();
 FILLCELL_X4 FILLER_0_85_793 ();
 FILLCELL_X1 FILLER_0_85_810 ();
 FILLCELL_X2 FILLER_0_85_818 ();
 FILLCELL_X1 FILLER_0_85_824 ();
 FILLCELL_X4 FILLER_0_85_842 ();
 FILLCELL_X2 FILLER_0_85_856 ();
 FILLCELL_X2 FILLER_0_85_868 ();
 FILLCELL_X4 FILLER_0_85_917 ();
 FILLCELL_X2 FILLER_0_85_938 ();
 FILLCELL_X1 FILLER_0_85_940 ();
 FILLCELL_X2 FILLER_0_85_958 ();
 FILLCELL_X1 FILLER_0_85_960 ();
 FILLCELL_X2 FILLER_0_85_983 ();
 FILLCELL_X1 FILLER_0_85_985 ();
 FILLCELL_X2 FILLER_0_85_996 ();
 FILLCELL_X4 FILLER_0_85_1013 ();
 FILLCELL_X1 FILLER_0_85_1022 ();
 FILLCELL_X8 FILLER_0_85_1033 ();
 FILLCELL_X4 FILLER_0_85_1041 ();
 FILLCELL_X2 FILLER_0_85_1045 ();
 FILLCELL_X2 FILLER_0_85_1126 ();
 FILLCELL_X32 FILLER_0_86_1 ();
 FILLCELL_X32 FILLER_0_86_33 ();
 FILLCELL_X32 FILLER_0_86_65 ();
 FILLCELL_X32 FILLER_0_86_97 ();
 FILLCELL_X32 FILLER_0_86_129 ();
 FILLCELL_X8 FILLER_0_86_161 ();
 FILLCELL_X4 FILLER_0_86_169 ();
 FILLCELL_X1 FILLER_0_86_173 ();
 FILLCELL_X2 FILLER_0_86_189 ();
 FILLCELL_X1 FILLER_0_86_191 ();
 FILLCELL_X2 FILLER_0_86_201 ();
 FILLCELL_X1 FILLER_0_86_203 ();
 FILLCELL_X8 FILLER_0_86_229 ();
 FILLCELL_X4 FILLER_0_86_237 ();
 FILLCELL_X2 FILLER_0_86_241 ();
 FILLCELL_X1 FILLER_0_86_243 ();
 FILLCELL_X1 FILLER_0_86_249 ();
 FILLCELL_X1 FILLER_0_86_320 ();
 FILLCELL_X2 FILLER_0_86_338 ();
 FILLCELL_X8 FILLER_0_86_370 ();
 FILLCELL_X2 FILLER_0_86_378 ();
 FILLCELL_X1 FILLER_0_86_380 ();
 FILLCELL_X8 FILLER_0_86_384 ();
 FILLCELL_X4 FILLER_0_86_392 ();
 FILLCELL_X2 FILLER_0_86_412 ();
 FILLCELL_X4 FILLER_0_86_468 ();
 FILLCELL_X2 FILLER_0_86_472 ();
 FILLCELL_X1 FILLER_0_86_474 ();
 FILLCELL_X1 FILLER_0_86_489 ();
 FILLCELL_X8 FILLER_0_86_493 ();
 FILLCELL_X1 FILLER_0_86_501 ();
 FILLCELL_X32 FILLER_0_86_524 ();
 FILLCELL_X8 FILLER_0_86_556 ();
 FILLCELL_X4 FILLER_0_86_564 ();
 FILLCELL_X8 FILLER_0_86_571 ();
 FILLCELL_X1 FILLER_0_86_579 ();
 FILLCELL_X8 FILLER_0_86_583 ();
 FILLCELL_X2 FILLER_0_86_591 ();
 FILLCELL_X1 FILLER_0_86_593 ();
 FILLCELL_X4 FILLER_0_86_624 ();
 FILLCELL_X2 FILLER_0_86_628 ();
 FILLCELL_X1 FILLER_0_86_630 ();
 FILLCELL_X1 FILLER_0_86_642 ();
 FILLCELL_X1 FILLER_0_86_653 ();
 FILLCELL_X1 FILLER_0_86_664 ();
 FILLCELL_X1 FILLER_0_86_670 ();
 FILLCELL_X16 FILLER_0_86_681 ();
 FILLCELL_X8 FILLER_0_86_697 ();
 FILLCELL_X4 FILLER_0_86_705 ();
 FILLCELL_X4 FILLER_0_86_719 ();
 FILLCELL_X1 FILLER_0_86_723 ();
 FILLCELL_X1 FILLER_0_86_739 ();
 FILLCELL_X2 FILLER_0_86_758 ();
 FILLCELL_X1 FILLER_0_86_760 ();
 FILLCELL_X4 FILLER_0_86_778 ();
 FILLCELL_X2 FILLER_0_86_782 ();
 FILLCELL_X1 FILLER_0_86_784 ();
 FILLCELL_X2 FILLER_0_86_798 ();
 FILLCELL_X2 FILLER_0_86_811 ();
 FILLCELL_X2 FILLER_0_86_823 ();
 FILLCELL_X1 FILLER_0_86_835 ();
 FILLCELL_X16 FILLER_0_86_850 ();
 FILLCELL_X4 FILLER_0_86_866 ();
 FILLCELL_X2 FILLER_0_86_870 ();
 FILLCELL_X4 FILLER_0_86_877 ();
 FILLCELL_X2 FILLER_0_86_881 ();
 FILLCELL_X1 FILLER_0_86_883 ();
 FILLCELL_X1 FILLER_0_86_889 ();
 FILLCELL_X2 FILLER_0_86_915 ();
 FILLCELL_X1 FILLER_0_86_917 ();
 FILLCELL_X4 FILLER_0_86_1003 ();
 FILLCELL_X1 FILLER_0_86_1007 ();
 FILLCELL_X8 FILLER_0_86_1038 ();
 FILLCELL_X4 FILLER_0_86_1046 ();
 FILLCELL_X1 FILLER_0_86_1050 ();
 FILLCELL_X1 FILLER_0_86_1058 ();
 FILLCELL_X4 FILLER_0_86_1090 ();
 FILLCELL_X2 FILLER_0_86_1146 ();
 FILLCELL_X32 FILLER_0_87_1 ();
 FILLCELL_X32 FILLER_0_87_33 ();
 FILLCELL_X32 FILLER_0_87_65 ();
 FILLCELL_X32 FILLER_0_87_97 ();
 FILLCELL_X32 FILLER_0_87_129 ();
 FILLCELL_X8 FILLER_0_87_161 ();
 FILLCELL_X4 FILLER_0_87_194 ();
 FILLCELL_X1 FILLER_0_87_198 ();
 FILLCELL_X4 FILLER_0_87_228 ();
 FILLCELL_X2 FILLER_0_87_232 ();
 FILLCELL_X1 FILLER_0_87_234 ();
 FILLCELL_X2 FILLER_0_87_245 ();
 FILLCELL_X4 FILLER_0_87_273 ();
 FILLCELL_X2 FILLER_0_87_292 ();
 FILLCELL_X1 FILLER_0_87_294 ();
 FILLCELL_X1 FILLER_0_87_335 ();
 FILLCELL_X8 FILLER_0_87_342 ();
 FILLCELL_X4 FILLER_0_87_350 ();
 FILLCELL_X2 FILLER_0_87_354 ();
 FILLCELL_X4 FILLER_0_87_360 ();
 FILLCELL_X1 FILLER_0_87_374 ();
 FILLCELL_X1 FILLER_0_87_379 ();
 FILLCELL_X2 FILLER_0_87_401 ();
 FILLCELL_X1 FILLER_0_87_403 ();
 FILLCELL_X2 FILLER_0_87_418 ();
 FILLCELL_X4 FILLER_0_87_423 ();
 FILLCELL_X1 FILLER_0_87_427 ();
 FILLCELL_X1 FILLER_0_87_453 ();
 FILLCELL_X8 FILLER_0_87_461 ();
 FILLCELL_X4 FILLER_0_87_469 ();
 FILLCELL_X4 FILLER_0_87_482 ();
 FILLCELL_X1 FILLER_0_87_486 ();
 FILLCELL_X1 FILLER_0_87_521 ();
 FILLCELL_X1 FILLER_0_87_524 ();
 FILLCELL_X1 FILLER_0_87_541 ();
 FILLCELL_X16 FILLER_0_87_551 ();
 FILLCELL_X1 FILLER_0_87_567 ();
 FILLCELL_X2 FILLER_0_87_578 ();
 FILLCELL_X8 FILLER_0_87_594 ();
 FILLCELL_X4 FILLER_0_87_602 ();
 FILLCELL_X2 FILLER_0_87_606 ();
 FILLCELL_X1 FILLER_0_87_608 ();
 FILLCELL_X2 FILLER_0_87_614 ();
 FILLCELL_X1 FILLER_0_87_616 ();
 FILLCELL_X2 FILLER_0_87_634 ();
 FILLCELL_X1 FILLER_0_87_636 ();
 FILLCELL_X2 FILLER_0_87_652 ();
 FILLCELL_X1 FILLER_0_87_654 ();
 FILLCELL_X4 FILLER_0_87_659 ();
 FILLCELL_X2 FILLER_0_87_663 ();
 FILLCELL_X1 FILLER_0_87_665 ();
 FILLCELL_X8 FILLER_0_87_670 ();
 FILLCELL_X4 FILLER_0_87_678 ();
 FILLCELL_X2 FILLER_0_87_682 ();
 FILLCELL_X4 FILLER_0_87_701 ();
 FILLCELL_X2 FILLER_0_87_705 ();
 FILLCELL_X1 FILLER_0_87_710 ();
 FILLCELL_X2 FILLER_0_87_716 ();
 FILLCELL_X1 FILLER_0_87_718 ();
 FILLCELL_X2 FILLER_0_87_729 ();
 FILLCELL_X2 FILLER_0_87_746 ();
 FILLCELL_X1 FILLER_0_87_761 ();
 FILLCELL_X2 FILLER_0_87_772 ();
 FILLCELL_X1 FILLER_0_87_774 ();
 FILLCELL_X2 FILLER_0_87_785 ();
 FILLCELL_X4 FILLER_0_87_860 ();
 FILLCELL_X1 FILLER_0_87_864 ();
 FILLCELL_X2 FILLER_0_87_886 ();
 FILLCELL_X1 FILLER_0_87_929 ();
 FILLCELL_X2 FILLER_0_87_935 ();
 FILLCELL_X2 FILLER_0_87_954 ();
 FILLCELL_X1 FILLER_0_87_956 ();
 FILLCELL_X4 FILLER_0_87_967 ();
 FILLCELL_X2 FILLER_0_87_981 ();
 FILLCELL_X8 FILLER_0_87_992 ();
 FILLCELL_X4 FILLER_0_87_1000 ();
 FILLCELL_X1 FILLER_0_87_1004 ();
 FILLCELL_X4 FILLER_0_87_1020 ();
 FILLCELL_X2 FILLER_0_87_1024 ();
 FILLCELL_X1 FILLER_0_87_1026 ();
 FILLCELL_X8 FILLER_0_87_1032 ();
 FILLCELL_X1 FILLER_0_87_1040 ();
 FILLCELL_X1 FILLER_0_87_1092 ();
 FILLCELL_X2 FILLER_0_87_1114 ();
 FILLCELL_X4 FILLER_0_87_1119 ();
 FILLCELL_X1 FILLER_0_87_1123 ();
 FILLCELL_X32 FILLER_0_88_1 ();
 FILLCELL_X32 FILLER_0_88_33 ();
 FILLCELL_X32 FILLER_0_88_65 ();
 FILLCELL_X32 FILLER_0_88_97 ();
 FILLCELL_X32 FILLER_0_88_129 ();
 FILLCELL_X16 FILLER_0_88_161 ();
 FILLCELL_X8 FILLER_0_88_177 ();
 FILLCELL_X4 FILLER_0_88_185 ();
 FILLCELL_X2 FILLER_0_88_189 ();
 FILLCELL_X2 FILLER_0_88_201 ();
 FILLCELL_X2 FILLER_0_88_222 ();
 FILLCELL_X1 FILLER_0_88_239 ();
 FILLCELL_X1 FILLER_0_88_250 ();
 FILLCELL_X2 FILLER_0_88_258 ();
 FILLCELL_X2 FILLER_0_88_270 ();
 FILLCELL_X8 FILLER_0_88_297 ();
 FILLCELL_X4 FILLER_0_88_310 ();
 FILLCELL_X2 FILLER_0_88_314 ();
 FILLCELL_X2 FILLER_0_88_326 ();
 FILLCELL_X1 FILLER_0_88_328 ();
 FILLCELL_X4 FILLER_0_88_346 ();
 FILLCELL_X2 FILLER_0_88_371 ();
 FILLCELL_X2 FILLER_0_88_414 ();
 FILLCELL_X1 FILLER_0_88_430 ();
 FILLCELL_X1 FILLER_0_88_438 ();
 FILLCELL_X2 FILLER_0_88_449 ();
 FILLCELL_X16 FILLER_0_88_454 ();
 FILLCELL_X1 FILLER_0_88_487 ();
 FILLCELL_X1 FILLER_0_88_498 ();
 FILLCELL_X4 FILLER_0_88_514 ();
 FILLCELL_X8 FILLER_0_88_553 ();
 FILLCELL_X2 FILLER_0_88_575 ();
 FILLCELL_X1 FILLER_0_88_577 ();
 FILLCELL_X1 FILLER_0_88_599 ();
 FILLCELL_X8 FILLER_0_88_603 ();
 FILLCELL_X1 FILLER_0_88_611 ();
 FILLCELL_X2 FILLER_0_88_629 ();
 FILLCELL_X4 FILLER_0_88_635 ();
 FILLCELL_X2 FILLER_0_88_639 ();
 FILLCELL_X1 FILLER_0_88_641 ();
 FILLCELL_X2 FILLER_0_88_678 ();
 FILLCELL_X1 FILLER_0_88_680 ();
 FILLCELL_X1 FILLER_0_88_696 ();
 FILLCELL_X1 FILLER_0_88_707 ();
 FILLCELL_X2 FILLER_0_88_712 ();
 FILLCELL_X2 FILLER_0_88_719 ();
 FILLCELL_X1 FILLER_0_88_721 ();
 FILLCELL_X1 FILLER_0_88_732 ();
 FILLCELL_X1 FILLER_0_88_753 ();
 FILLCELL_X4 FILLER_0_88_764 ();
 FILLCELL_X1 FILLER_0_88_768 ();
 FILLCELL_X2 FILLER_0_88_773 ();
 FILLCELL_X1 FILLER_0_88_775 ();
 FILLCELL_X2 FILLER_0_88_895 ();
 FILLCELL_X2 FILLER_0_88_946 ();
 FILLCELL_X2 FILLER_0_88_973 ();
 FILLCELL_X1 FILLER_0_88_985 ();
 FILLCELL_X4 FILLER_0_88_991 ();
 FILLCELL_X2 FILLER_0_88_995 ();
 FILLCELL_X1 FILLER_0_88_997 ();
 FILLCELL_X2 FILLER_0_88_1008 ();
 FILLCELL_X8 FILLER_0_88_1035 ();
 FILLCELL_X1 FILLER_0_88_1140 ();
 FILLCELL_X32 FILLER_0_89_1 ();
 FILLCELL_X32 FILLER_0_89_33 ();
 FILLCELL_X32 FILLER_0_89_65 ();
 FILLCELL_X32 FILLER_0_89_97 ();
 FILLCELL_X32 FILLER_0_89_129 ();
 FILLCELL_X32 FILLER_0_89_161 ();
 FILLCELL_X2 FILLER_0_89_193 ();
 FILLCELL_X1 FILLER_0_89_195 ();
 FILLCELL_X1 FILLER_0_89_206 ();
 FILLCELL_X1 FILLER_0_89_212 ();
 FILLCELL_X1 FILLER_0_89_218 ();
 FILLCELL_X1 FILLER_0_89_226 ();
 FILLCELL_X8 FILLER_0_89_237 ();
 FILLCELL_X2 FILLER_0_89_245 ();
 FILLCELL_X32 FILLER_0_89_254 ();
 FILLCELL_X16 FILLER_0_89_293 ();
 FILLCELL_X8 FILLER_0_89_309 ();
 FILLCELL_X2 FILLER_0_89_317 ();
 FILLCELL_X1 FILLER_0_89_319 ();
 FILLCELL_X4 FILLER_0_89_351 ();
 FILLCELL_X2 FILLER_0_89_355 ();
 FILLCELL_X8 FILLER_0_89_362 ();
 FILLCELL_X2 FILLER_0_89_370 ();
 FILLCELL_X1 FILLER_0_89_372 ();
 FILLCELL_X1 FILLER_0_89_395 ();
 FILLCELL_X4 FILLER_0_89_411 ();
 FILLCELL_X4 FILLER_0_89_430 ();
 FILLCELL_X1 FILLER_0_89_434 ();
 FILLCELL_X4 FILLER_0_89_466 ();
 FILLCELL_X8 FILLER_0_89_473 ();
 FILLCELL_X4 FILLER_0_89_481 ();
 FILLCELL_X1 FILLER_0_89_485 ();
 FILLCELL_X2 FILLER_0_89_542 ();
 FILLCELL_X4 FILLER_0_89_561 ();
 FILLCELL_X1 FILLER_0_89_565 ();
 FILLCELL_X8 FILLER_0_89_588 ();
 FILLCELL_X4 FILLER_0_89_596 ();
 FILLCELL_X2 FILLER_0_89_614 ();
 FILLCELL_X1 FILLER_0_89_616 ();
 FILLCELL_X2 FILLER_0_89_648 ();
 FILLCELL_X1 FILLER_0_89_650 ();
 FILLCELL_X1 FILLER_0_89_668 ();
 FILLCELL_X1 FILLER_0_89_683 ();
 FILLCELL_X2 FILLER_0_89_701 ();
 FILLCELL_X1 FILLER_0_89_703 ();
 FILLCELL_X2 FILLER_0_89_724 ();
 FILLCELL_X8 FILLER_0_89_740 ();
 FILLCELL_X1 FILLER_0_89_748 ();
 FILLCELL_X8 FILLER_0_89_759 ();
 FILLCELL_X2 FILLER_0_89_767 ();
 FILLCELL_X1 FILLER_0_89_769 ();
 FILLCELL_X1 FILLER_0_89_836 ();
 FILLCELL_X4 FILLER_0_89_898 ();
 FILLCELL_X1 FILLER_0_89_902 ();
 FILLCELL_X4 FILLER_0_89_913 ();
 FILLCELL_X1 FILLER_0_89_917 ();
 FILLCELL_X2 FILLER_0_89_991 ();
 FILLCELL_X8 FILLER_0_89_1023 ();
 FILLCELL_X4 FILLER_0_89_1031 ();
 FILLCELL_X1 FILLER_0_89_1035 ();
 FILLCELL_X1 FILLER_0_89_1147 ();
 FILLCELL_X32 FILLER_0_90_1 ();
 FILLCELL_X32 FILLER_0_90_33 ();
 FILLCELL_X32 FILLER_0_90_65 ();
 FILLCELL_X32 FILLER_0_90_97 ();
 FILLCELL_X32 FILLER_0_90_129 ();
 FILLCELL_X32 FILLER_0_90_161 ();
 FILLCELL_X8 FILLER_0_90_193 ();
 FILLCELL_X4 FILLER_0_90_201 ();
 FILLCELL_X2 FILLER_0_90_205 ();
 FILLCELL_X1 FILLER_0_90_207 ();
 FILLCELL_X32 FILLER_0_90_218 ();
 FILLCELL_X4 FILLER_0_90_250 ();
 FILLCELL_X4 FILLER_0_90_264 ();
 FILLCELL_X1 FILLER_0_90_268 ();
 FILLCELL_X1 FILLER_0_90_289 ();
 FILLCELL_X2 FILLER_0_90_324 ();
 FILLCELL_X4 FILLER_0_90_346 ();
 FILLCELL_X1 FILLER_0_90_370 ();
 FILLCELL_X1 FILLER_0_90_391 ();
 FILLCELL_X1 FILLER_0_90_403 ();
 FILLCELL_X8 FILLER_0_90_414 ();
 FILLCELL_X1 FILLER_0_90_422 ();
 FILLCELL_X1 FILLER_0_90_447 ();
 FILLCELL_X2 FILLER_0_90_468 ();
 FILLCELL_X1 FILLER_0_90_480 ();
 FILLCELL_X2 FILLER_0_90_502 ();
 FILLCELL_X4 FILLER_0_90_543 ();
 FILLCELL_X2 FILLER_0_90_547 ();
 FILLCELL_X1 FILLER_0_90_549 ();
 FILLCELL_X1 FILLER_0_90_560 ();
 FILLCELL_X4 FILLER_0_90_571 ();
 FILLCELL_X4 FILLER_0_90_600 ();
 FILLCELL_X2 FILLER_0_90_604 ();
 FILLCELL_X1 FILLER_0_90_609 ();
 FILLCELL_X2 FILLER_0_90_620 ();
 FILLCELL_X2 FILLER_0_90_629 ();
 FILLCELL_X1 FILLER_0_90_635 ();
 FILLCELL_X2 FILLER_0_90_652 ();
 FILLCELL_X1 FILLER_0_90_667 ();
 FILLCELL_X2 FILLER_0_90_675 ();
 FILLCELL_X1 FILLER_0_90_709 ();
 FILLCELL_X1 FILLER_0_90_713 ();
 FILLCELL_X2 FILLER_0_90_754 ();
 FILLCELL_X2 FILLER_0_90_766 ();
 FILLCELL_X1 FILLER_0_90_768 ();
 FILLCELL_X2 FILLER_0_90_774 ();
 FILLCELL_X1 FILLER_0_90_776 ();
 FILLCELL_X2 FILLER_0_90_786 ();
 FILLCELL_X2 FILLER_0_90_822 ();
 FILLCELL_X1 FILLER_0_90_847 ();
 FILLCELL_X1 FILLER_0_90_867 ();
 FILLCELL_X1 FILLER_0_90_875 ();
 FILLCELL_X1 FILLER_0_90_879 ();
 FILLCELL_X16 FILLER_0_90_901 ();
 FILLCELL_X4 FILLER_0_90_917 ();
 FILLCELL_X1 FILLER_0_90_921 ();
 FILLCELL_X2 FILLER_0_90_937 ();
 FILLCELL_X16 FILLER_0_90_953 ();
 FILLCELL_X4 FILLER_0_90_969 ();
 FILLCELL_X2 FILLER_0_90_973 ();
 FILLCELL_X1 FILLER_0_90_1000 ();
 FILLCELL_X2 FILLER_0_90_1006 ();
 FILLCELL_X1 FILLER_0_90_1008 ();
 FILLCELL_X16 FILLER_0_90_1014 ();
 FILLCELL_X8 FILLER_0_90_1030 ();
 FILLCELL_X32 FILLER_0_91_1 ();
 FILLCELL_X32 FILLER_0_91_33 ();
 FILLCELL_X32 FILLER_0_91_65 ();
 FILLCELL_X32 FILLER_0_91_97 ();
 FILLCELL_X32 FILLER_0_91_129 ();
 FILLCELL_X32 FILLER_0_91_161 ();
 FILLCELL_X32 FILLER_0_91_193 ();
 FILLCELL_X16 FILLER_0_91_225 ();
 FILLCELL_X8 FILLER_0_91_241 ();
 FILLCELL_X2 FILLER_0_91_249 ();
 FILLCELL_X1 FILLER_0_91_251 ();
 FILLCELL_X2 FILLER_0_91_269 ();
 FILLCELL_X1 FILLER_0_91_276 ();
 FILLCELL_X2 FILLER_0_91_287 ();
 FILLCELL_X4 FILLER_0_91_324 ();
 FILLCELL_X1 FILLER_0_91_328 ();
 FILLCELL_X8 FILLER_0_91_333 ();
 FILLCELL_X4 FILLER_0_91_341 ();
 FILLCELL_X4 FILLER_0_91_348 ();
 FILLCELL_X2 FILLER_0_91_352 ();
 FILLCELL_X1 FILLER_0_91_354 ();
 FILLCELL_X2 FILLER_0_91_368 ();
 FILLCELL_X2 FILLER_0_91_374 ();
 FILLCELL_X4 FILLER_0_91_427 ();
 FILLCELL_X1 FILLER_0_91_431 ();
 FILLCELL_X2 FILLER_0_91_436 ();
 FILLCELL_X4 FILLER_0_91_471 ();
 FILLCELL_X1 FILLER_0_91_475 ();
 FILLCELL_X4 FILLER_0_91_486 ();
 FILLCELL_X2 FILLER_0_91_490 ();
 FILLCELL_X4 FILLER_0_91_516 ();
 FILLCELL_X2 FILLER_0_91_520 ();
 FILLCELL_X1 FILLER_0_91_532 ();
 FILLCELL_X4 FILLER_0_91_550 ();
 FILLCELL_X8 FILLER_0_91_607 ();
 FILLCELL_X2 FILLER_0_91_615 ();
 FILLCELL_X1 FILLER_0_91_617 ();
 FILLCELL_X4 FILLER_0_91_622 ();
 FILLCELL_X1 FILLER_0_91_626 ();
 FILLCELL_X4 FILLER_0_91_662 ();
 FILLCELL_X1 FILLER_0_91_676 ();
 FILLCELL_X2 FILLER_0_91_691 ();
 FILLCELL_X1 FILLER_0_91_708 ();
 FILLCELL_X2 FILLER_0_91_745 ();
 FILLCELL_X8 FILLER_0_91_757 ();
 FILLCELL_X1 FILLER_0_91_792 ();
 FILLCELL_X1 FILLER_0_91_846 ();
 FILLCELL_X2 FILLER_0_91_857 ();
 FILLCELL_X1 FILLER_0_91_859 ();
 FILLCELL_X1 FILLER_0_91_863 ();
 FILLCELL_X16 FILLER_0_91_909 ();
 FILLCELL_X8 FILLER_0_91_925 ();
 FILLCELL_X1 FILLER_0_91_933 ();
 FILLCELL_X32 FILLER_0_91_964 ();
 FILLCELL_X4 FILLER_0_91_996 ();
 FILLCELL_X2 FILLER_0_91_1000 ();
 FILLCELL_X16 FILLER_0_91_1012 ();
 FILLCELL_X4 FILLER_0_91_1028 ();
 FILLCELL_X2 FILLER_0_91_1032 ();
 FILLCELL_X1 FILLER_0_91_1034 ();
 FILLCELL_X2 FILLER_0_91_1081 ();
 FILLCELL_X32 FILLER_0_92_1 ();
 FILLCELL_X32 FILLER_0_92_33 ();
 FILLCELL_X32 FILLER_0_92_65 ();
 FILLCELL_X32 FILLER_0_92_97 ();
 FILLCELL_X32 FILLER_0_92_129 ();
 FILLCELL_X32 FILLER_0_92_161 ();
 FILLCELL_X16 FILLER_0_92_193 ();
 FILLCELL_X8 FILLER_0_92_209 ();
 FILLCELL_X1 FILLER_0_92_227 ();
 FILLCELL_X4 FILLER_0_92_238 ();
 FILLCELL_X1 FILLER_0_92_242 ();
 FILLCELL_X8 FILLER_0_92_247 ();
 FILLCELL_X1 FILLER_0_92_265 ();
 FILLCELL_X1 FILLER_0_92_276 ();
 FILLCELL_X1 FILLER_0_92_282 ();
 FILLCELL_X2 FILLER_0_92_339 ();
 FILLCELL_X2 FILLER_0_92_355 ();
 FILLCELL_X1 FILLER_0_92_375 ();
 FILLCELL_X1 FILLER_0_92_406 ();
 FILLCELL_X2 FILLER_0_92_421 ();
 FILLCELL_X1 FILLER_0_92_430 ();
 FILLCELL_X8 FILLER_0_92_438 ();
 FILLCELL_X1 FILLER_0_92_467 ();
 FILLCELL_X2 FILLER_0_92_482 ();
 FILLCELL_X1 FILLER_0_92_517 ();
 FILLCELL_X4 FILLER_0_92_528 ();
 FILLCELL_X1 FILLER_0_92_532 ();
 FILLCELL_X2 FILLER_0_92_555 ();
 FILLCELL_X2 FILLER_0_92_562 ();
 FILLCELL_X1 FILLER_0_92_564 ();
 FILLCELL_X2 FILLER_0_92_574 ();
 FILLCELL_X4 FILLER_0_92_606 ();
 FILLCELL_X2 FILLER_0_92_610 ();
 FILLCELL_X2 FILLER_0_92_626 ();
 FILLCELL_X2 FILLER_0_92_632 ();
 FILLCELL_X1 FILLER_0_92_659 ();
 FILLCELL_X2 FILLER_0_92_670 ();
 FILLCELL_X2 FILLER_0_92_686 ();
 FILLCELL_X2 FILLER_0_92_741 ();
 FILLCELL_X4 FILLER_0_92_754 ();
 FILLCELL_X2 FILLER_0_92_758 ();
 FILLCELL_X1 FILLER_0_92_760 ();
 FILLCELL_X2 FILLER_0_92_766 ();
 FILLCELL_X1 FILLER_0_92_768 ();
 FILLCELL_X8 FILLER_0_92_812 ();
 FILLCELL_X4 FILLER_0_92_820 ();
 FILLCELL_X2 FILLER_0_92_824 ();
 FILLCELL_X2 FILLER_0_92_846 ();
 FILLCELL_X1 FILLER_0_92_858 ();
 FILLCELL_X1 FILLER_0_92_870 ();
 FILLCELL_X4 FILLER_0_92_916 ();
 FILLCELL_X2 FILLER_0_92_920 ();
 FILLCELL_X4 FILLER_0_92_947 ();
 FILLCELL_X1 FILLER_0_92_961 ();
 FILLCELL_X4 FILLER_0_92_972 ();
 FILLCELL_X1 FILLER_0_92_976 ();
 FILLCELL_X2 FILLER_0_92_987 ();
 FILLCELL_X16 FILLER_0_92_998 ();
 FILLCELL_X8 FILLER_0_92_1014 ();
 FILLCELL_X4 FILLER_0_92_1022 ();
 FILLCELL_X32 FILLER_0_93_1 ();
 FILLCELL_X32 FILLER_0_93_33 ();
 FILLCELL_X32 FILLER_0_93_65 ();
 FILLCELL_X32 FILLER_0_93_97 ();
 FILLCELL_X32 FILLER_0_93_129 ();
 FILLCELL_X32 FILLER_0_93_161 ();
 FILLCELL_X8 FILLER_0_93_193 ();
 FILLCELL_X4 FILLER_0_93_201 ();
 FILLCELL_X1 FILLER_0_93_205 ();
 FILLCELL_X1 FILLER_0_93_221 ();
 FILLCELL_X1 FILLER_0_93_236 ();
 FILLCELL_X1 FILLER_0_93_266 ();
 FILLCELL_X1 FILLER_0_93_305 ();
 FILLCELL_X2 FILLER_0_93_308 ();
 FILLCELL_X1 FILLER_0_93_320 ();
 FILLCELL_X1 FILLER_0_93_331 ();
 FILLCELL_X2 FILLER_0_93_347 ();
 FILLCELL_X1 FILLER_0_93_349 ();
 FILLCELL_X2 FILLER_0_93_360 ();
 FILLCELL_X1 FILLER_0_93_407 ();
 FILLCELL_X2 FILLER_0_93_447 ();
 FILLCELL_X8 FILLER_0_93_467 ();
 FILLCELL_X2 FILLER_0_93_475 ();
 FILLCELL_X1 FILLER_0_93_477 ();
 FILLCELL_X4 FILLER_0_93_516 ();
 FILLCELL_X1 FILLER_0_93_566 ();
 FILLCELL_X8 FILLER_0_93_592 ();
 FILLCELL_X2 FILLER_0_93_600 ();
 FILLCELL_X1 FILLER_0_93_602 ();
 FILLCELL_X2 FILLER_0_93_613 ();
 FILLCELL_X8 FILLER_0_93_636 ();
 FILLCELL_X4 FILLER_0_93_644 ();
 FILLCELL_X2 FILLER_0_93_648 ();
 FILLCELL_X1 FILLER_0_93_681 ();
 FILLCELL_X2 FILLER_0_93_785 ();
 FILLCELL_X2 FILLER_0_93_797 ();
 FILLCELL_X1 FILLER_0_93_799 ();
 FILLCELL_X8 FILLER_0_93_820 ();
 FILLCELL_X2 FILLER_0_93_828 ();
 FILLCELL_X2 FILLER_0_93_850 ();
 FILLCELL_X1 FILLER_0_93_862 ();
 FILLCELL_X1 FILLER_0_93_898 ();
 FILLCELL_X2 FILLER_0_93_903 ();
 FILLCELL_X1 FILLER_0_93_905 ();
 FILLCELL_X4 FILLER_0_93_921 ();
 FILLCELL_X2 FILLER_0_93_925 ();
 FILLCELL_X1 FILLER_0_93_927 ();
 FILLCELL_X4 FILLER_0_93_942 ();
 FILLCELL_X2 FILLER_0_93_946 ();
 FILLCELL_X1 FILLER_0_93_963 ();
 FILLCELL_X4 FILLER_0_93_1006 ();
 FILLCELL_X2 FILLER_0_93_1010 ();
 FILLCELL_X1 FILLER_0_93_1012 ();
 FILLCELL_X4 FILLER_0_93_1023 ();
 FILLCELL_X1 FILLER_0_93_1027 ();
 FILLCELL_X2 FILLER_0_93_1033 ();
 FILLCELL_X4 FILLER_0_93_1045 ();
 FILLCELL_X2 FILLER_0_93_1049 ();
 FILLCELL_X1 FILLER_0_93_1051 ();
 FILLCELL_X1 FILLER_0_93_1111 ();
 FILLCELL_X2 FILLER_0_93_1139 ();
 FILLCELL_X32 FILLER_0_94_1 ();
 FILLCELL_X32 FILLER_0_94_33 ();
 FILLCELL_X32 FILLER_0_94_65 ();
 FILLCELL_X32 FILLER_0_94_97 ();
 FILLCELL_X32 FILLER_0_94_129 ();
 FILLCELL_X32 FILLER_0_94_161 ();
 FILLCELL_X16 FILLER_0_94_193 ();
 FILLCELL_X4 FILLER_0_94_209 ();
 FILLCELL_X1 FILLER_0_94_213 ();
 FILLCELL_X2 FILLER_0_94_234 ();
 FILLCELL_X1 FILLER_0_94_236 ();
 FILLCELL_X1 FILLER_0_94_247 ();
 FILLCELL_X2 FILLER_0_94_297 ();
 FILLCELL_X4 FILLER_0_94_305 ();
 FILLCELL_X1 FILLER_0_94_320 ();
 FILLCELL_X2 FILLER_0_94_335 ();
 FILLCELL_X2 FILLER_0_94_358 ();
 FILLCELL_X1 FILLER_0_94_384 ();
 FILLCELL_X1 FILLER_0_94_445 ();
 FILLCELL_X1 FILLER_0_94_466 ();
 FILLCELL_X2 FILLER_0_94_470 ();
 FILLCELL_X1 FILLER_0_94_472 ();
 FILLCELL_X2 FILLER_0_94_485 ();
 FILLCELL_X1 FILLER_0_94_487 ();
 FILLCELL_X2 FILLER_0_94_493 ();
 FILLCELL_X1 FILLER_0_94_495 ();
 FILLCELL_X1 FILLER_0_94_539 ();
 FILLCELL_X2 FILLER_0_94_555 ();
 FILLCELL_X4 FILLER_0_94_567 ();
 FILLCELL_X1 FILLER_0_94_571 ();
 FILLCELL_X2 FILLER_0_94_577 ();
 FILLCELL_X8 FILLER_0_94_589 ();
 FILLCELL_X2 FILLER_0_94_629 ();
 FILLCELL_X4 FILLER_0_94_635 ();
 FILLCELL_X2 FILLER_0_94_639 ();
 FILLCELL_X4 FILLER_0_94_659 ();
 FILLCELL_X2 FILLER_0_94_663 ();
 FILLCELL_X1 FILLER_0_94_688 ();
 FILLCELL_X2 FILLER_0_94_730 ();
 FILLCELL_X2 FILLER_0_94_742 ();
 FILLCELL_X1 FILLER_0_94_754 ();
 FILLCELL_X1 FILLER_0_94_777 ();
 FILLCELL_X1 FILLER_0_94_793 ();
 FILLCELL_X2 FILLER_0_94_804 ();
 FILLCELL_X4 FILLER_0_94_823 ();
 FILLCELL_X2 FILLER_0_94_827 ();
 FILLCELL_X1 FILLER_0_94_829 ();
 FILLCELL_X2 FILLER_0_94_862 ();
 FILLCELL_X8 FILLER_0_94_896 ();
 FILLCELL_X4 FILLER_0_94_904 ();
 FILLCELL_X2 FILLER_0_94_908 ();
 FILLCELL_X1 FILLER_0_94_910 ();
 FILLCELL_X4 FILLER_0_94_915 ();
 FILLCELL_X8 FILLER_0_94_934 ();
 FILLCELL_X1 FILLER_0_94_942 ();
 FILLCELL_X1 FILLER_0_94_968 ();
 FILLCELL_X1 FILLER_0_94_1016 ();
 FILLCELL_X2 FILLER_0_94_1027 ();
 FILLCELL_X1 FILLER_0_94_1090 ();
 FILLCELL_X1 FILLER_0_94_1118 ();
 FILLCELL_X2 FILLER_0_94_1139 ();
 FILLCELL_X32 FILLER_0_95_1 ();
 FILLCELL_X32 FILLER_0_95_33 ();
 FILLCELL_X32 FILLER_0_95_65 ();
 FILLCELL_X32 FILLER_0_95_97 ();
 FILLCELL_X32 FILLER_0_95_129 ();
 FILLCELL_X32 FILLER_0_95_161 ();
 FILLCELL_X32 FILLER_0_95_193 ();
 FILLCELL_X1 FILLER_0_95_225 ();
 FILLCELL_X16 FILLER_0_95_236 ();
 FILLCELL_X1 FILLER_0_95_252 ();
 FILLCELL_X1 FILLER_0_95_263 ();
 FILLCELL_X2 FILLER_0_95_279 ();
 FILLCELL_X1 FILLER_0_95_281 ();
 FILLCELL_X4 FILLER_0_95_305 ();
 FILLCELL_X1 FILLER_0_95_328 ();
 FILLCELL_X1 FILLER_0_95_333 ();
 FILLCELL_X4 FILLER_0_95_347 ();
 FILLCELL_X1 FILLER_0_95_351 ();
 FILLCELL_X1 FILLER_0_95_407 ();
 FILLCELL_X1 FILLER_0_95_436 ();
 FILLCELL_X2 FILLER_0_95_447 ();
 FILLCELL_X1 FILLER_0_95_471 ();
 FILLCELL_X2 FILLER_0_95_482 ();
 FILLCELL_X1 FILLER_0_95_491 ();
 FILLCELL_X2 FILLER_0_95_503 ();
 FILLCELL_X2 FILLER_0_95_556 ();
 FILLCELL_X1 FILLER_0_95_573 ();
 FILLCELL_X1 FILLER_0_95_584 ();
 FILLCELL_X8 FILLER_0_95_595 ();
 FILLCELL_X1 FILLER_0_95_603 ();
 FILLCELL_X1 FILLER_0_95_624 ();
 FILLCELL_X1 FILLER_0_95_628 ();
 FILLCELL_X2 FILLER_0_95_643 ();
 FILLCELL_X2 FILLER_0_95_682 ();
 FILLCELL_X1 FILLER_0_95_684 ();
 FILLCELL_X2 FILLER_0_95_690 ();
 FILLCELL_X1 FILLER_0_95_702 ();
 FILLCELL_X2 FILLER_0_95_715 ();
 FILLCELL_X2 FILLER_0_95_748 ();
 FILLCELL_X1 FILLER_0_95_750 ();
 FILLCELL_X1 FILLER_0_95_811 ();
 FILLCELL_X2 FILLER_0_95_822 ();
 FILLCELL_X4 FILLER_0_95_831 ();
 FILLCELL_X1 FILLER_0_95_835 ();
 FILLCELL_X1 FILLER_0_95_853 ();
 FILLCELL_X1 FILLER_0_95_858 ();
 FILLCELL_X2 FILLER_0_95_863 ();
 FILLCELL_X2 FILLER_0_95_892 ();
 FILLCELL_X16 FILLER_0_95_904 ();
 FILLCELL_X2 FILLER_0_95_920 ();
 FILLCELL_X1 FILLER_0_95_947 ();
 FILLCELL_X2 FILLER_0_95_983 ();
 FILLCELL_X1 FILLER_0_95_985 ();
 FILLCELL_X4 FILLER_0_95_996 ();
 FILLCELL_X2 FILLER_0_95_1015 ();
 FILLCELL_X1 FILLER_0_95_1027 ();
 FILLCELL_X8 FILLER_0_95_1038 ();
 FILLCELL_X4 FILLER_0_95_1046 ();
 FILLCELL_X32 FILLER_0_96_1 ();
 FILLCELL_X32 FILLER_0_96_33 ();
 FILLCELL_X32 FILLER_0_96_65 ();
 FILLCELL_X32 FILLER_0_96_97 ();
 FILLCELL_X32 FILLER_0_96_129 ();
 FILLCELL_X32 FILLER_0_96_161 ();
 FILLCELL_X16 FILLER_0_96_193 ();
 FILLCELL_X8 FILLER_0_96_209 ();
 FILLCELL_X4 FILLER_0_96_217 ();
 FILLCELL_X1 FILLER_0_96_221 ();
 FILLCELL_X1 FILLER_0_96_247 ();
 FILLCELL_X2 FILLER_0_96_258 ();
 FILLCELL_X2 FILLER_0_96_297 ();
 FILLCELL_X1 FILLER_0_96_309 ();
 FILLCELL_X2 FILLER_0_96_427 ();
 FILLCELL_X4 FILLER_0_96_433 ();
 FILLCELL_X1 FILLER_0_96_437 ();
 FILLCELL_X1 FILLER_0_96_455 ();
 FILLCELL_X1 FILLER_0_96_466 ();
 FILLCELL_X2 FILLER_0_96_477 ();
 FILLCELL_X2 FILLER_0_96_483 ();
 FILLCELL_X1 FILLER_0_96_498 ();
 FILLCELL_X1 FILLER_0_96_562 ();
 FILLCELL_X2 FILLER_0_96_573 ();
 FILLCELL_X1 FILLER_0_96_575 ();
 FILLCELL_X2 FILLER_0_96_581 ();
 FILLCELL_X1 FILLER_0_96_583 ();
 FILLCELL_X1 FILLER_0_96_589 ();
 FILLCELL_X4 FILLER_0_96_669 ();
 FILLCELL_X2 FILLER_0_96_688 ();
 FILLCELL_X1 FILLER_0_96_690 ();
 FILLCELL_X1 FILLER_0_96_738 ();
 FILLCELL_X2 FILLER_0_96_775 ();
 FILLCELL_X1 FILLER_0_96_784 ();
 FILLCELL_X8 FILLER_0_96_820 ();
 FILLCELL_X1 FILLER_0_96_828 ();
 FILLCELL_X2 FILLER_0_96_856 ();
 FILLCELL_X1 FILLER_0_96_868 ();
 FILLCELL_X2 FILLER_0_96_929 ();
 FILLCELL_X1 FILLER_0_96_931 ();
 FILLCELL_X2 FILLER_0_96_957 ();
 FILLCELL_X2 FILLER_0_96_976 ();
 FILLCELL_X2 FILLER_0_96_1017 ();
 FILLCELL_X2 FILLER_0_96_1024 ();
 FILLCELL_X1 FILLER_0_96_1026 ();
 FILLCELL_X1 FILLER_0_96_1032 ();
 FILLCELL_X4 FILLER_0_96_1065 ();
 FILLCELL_X2 FILLER_0_96_1103 ();
 FILLCELL_X1 FILLER_0_96_1147 ();
 FILLCELL_X32 FILLER_0_97_1 ();
 FILLCELL_X32 FILLER_0_97_33 ();
 FILLCELL_X32 FILLER_0_97_65 ();
 FILLCELL_X32 FILLER_0_97_97 ();
 FILLCELL_X32 FILLER_0_97_129 ();
 FILLCELL_X32 FILLER_0_97_161 ();
 FILLCELL_X8 FILLER_0_97_193 ();
 FILLCELL_X4 FILLER_0_97_201 ();
 FILLCELL_X1 FILLER_0_97_205 ();
 FILLCELL_X2 FILLER_0_97_230 ();
 FILLCELL_X1 FILLER_0_97_232 ();
 FILLCELL_X2 FILLER_0_97_270 ();
 FILLCELL_X1 FILLER_0_97_272 ();
 FILLCELL_X2 FILLER_0_97_305 ();
 FILLCELL_X2 FILLER_0_97_412 ();
 FILLCELL_X4 FILLER_0_97_437 ();
 FILLCELL_X2 FILLER_0_97_441 ();
 FILLCELL_X1 FILLER_0_97_443 ();
 FILLCELL_X2 FILLER_0_97_484 ();
 FILLCELL_X2 FILLER_0_97_496 ();
 FILLCELL_X2 FILLER_0_97_519 ();
 FILLCELL_X1 FILLER_0_97_521 ();
 FILLCELL_X1 FILLER_0_97_532 ();
 FILLCELL_X2 FILLER_0_97_562 ();
 FILLCELL_X4 FILLER_0_97_574 ();
 FILLCELL_X4 FILLER_0_97_591 ();
 FILLCELL_X2 FILLER_0_97_600 ();
 FILLCELL_X2 FILLER_0_97_612 ();
 FILLCELL_X2 FILLER_0_97_624 ();
 FILLCELL_X1 FILLER_0_97_626 ();
 FILLCELL_X2 FILLER_0_97_650 ();
 FILLCELL_X4 FILLER_0_97_663 ();
 FILLCELL_X1 FILLER_0_97_667 ();
 FILLCELL_X1 FILLER_0_97_717 ();
 FILLCELL_X1 FILLER_0_97_725 ();
 FILLCELL_X1 FILLER_0_97_733 ();
 FILLCELL_X1 FILLER_0_97_749 ();
 FILLCELL_X2 FILLER_0_97_822 ();
 FILLCELL_X1 FILLER_0_97_824 ();
 FILLCELL_X1 FILLER_0_97_828 ();
 FILLCELL_X1 FILLER_0_97_925 ();
 FILLCELL_X2 FILLER_0_97_936 ();
 FILLCELL_X1 FILLER_0_97_938 ();
 FILLCELL_X2 FILLER_0_97_970 ();
 FILLCELL_X4 FILLER_0_97_1044 ();
 FILLCELL_X2 FILLER_0_97_1070 ();
 FILLCELL_X2 FILLER_0_97_1105 ();
 FILLCELL_X2 FILLER_0_97_1126 ();
 FILLCELL_X32 FILLER_0_98_1 ();
 FILLCELL_X32 FILLER_0_98_33 ();
 FILLCELL_X32 FILLER_0_98_65 ();
 FILLCELL_X32 FILLER_0_98_97 ();
 FILLCELL_X32 FILLER_0_98_129 ();
 FILLCELL_X32 FILLER_0_98_161 ();
 FILLCELL_X16 FILLER_0_98_193 ();
 FILLCELL_X2 FILLER_0_98_234 ();
 FILLCELL_X1 FILLER_0_98_236 ();
 FILLCELL_X1 FILLER_0_98_329 ();
 FILLCELL_X1 FILLER_0_98_385 ();
 FILLCELL_X4 FILLER_0_98_438 ();
 FILLCELL_X2 FILLER_0_98_442 ();
 FILLCELL_X2 FILLER_0_98_454 ();
 FILLCELL_X1 FILLER_0_98_456 ();
 FILLCELL_X1 FILLER_0_98_504 ();
 FILLCELL_X1 FILLER_0_98_541 ();
 FILLCELL_X1 FILLER_0_98_556 ();
 FILLCELL_X8 FILLER_0_98_589 ();
 FILLCELL_X16 FILLER_0_98_607 ();
 FILLCELL_X8 FILLER_0_98_623 ();
 FILLCELL_X1 FILLER_0_98_635 ();
 FILLCELL_X1 FILLER_0_98_646 ();
 FILLCELL_X1 FILLER_0_98_673 ();
 FILLCELL_X1 FILLER_0_98_752 ();
 FILLCELL_X4 FILLER_0_98_811 ();
 FILLCELL_X2 FILLER_0_98_823 ();
 FILLCELL_X1 FILLER_0_98_825 ();
 FILLCELL_X2 FILLER_0_98_836 ();
 FILLCELL_X1 FILLER_0_98_838 ();
 FILLCELL_X1 FILLER_0_98_862 ();
 FILLCELL_X2 FILLER_0_98_943 ();
 FILLCELL_X1 FILLER_0_98_945 ();
 FILLCELL_X2 FILLER_0_98_982 ();
 FILLCELL_X2 FILLER_0_98_1001 ();
 FILLCELL_X2 FILLER_0_98_1013 ();
 FILLCELL_X1 FILLER_0_98_1015 ();
 FILLCELL_X2 FILLER_0_98_1033 ();
 FILLCELL_X1 FILLER_0_98_1035 ();
 FILLCELL_X2 FILLER_0_98_1046 ();
 FILLCELL_X1 FILLER_0_98_1048 ();
 FILLCELL_X2 FILLER_0_98_1063 ();
 FILLCELL_X4 FILLER_0_98_1087 ();
 FILLCELL_X2 FILLER_0_98_1091 ();
 FILLCELL_X2 FILLER_0_98_1108 ();
 FILLCELL_X2 FILLER_0_98_1146 ();
 FILLCELL_X32 FILLER_0_99_1 ();
 FILLCELL_X32 FILLER_0_99_33 ();
 FILLCELL_X32 FILLER_0_99_65 ();
 FILLCELL_X32 FILLER_0_99_97 ();
 FILLCELL_X32 FILLER_0_99_129 ();
 FILLCELL_X32 FILLER_0_99_161 ();
 FILLCELL_X16 FILLER_0_99_193 ();
 FILLCELL_X8 FILLER_0_99_209 ();
 FILLCELL_X2 FILLER_0_99_217 ();
 FILLCELL_X2 FILLER_0_99_239 ();
 FILLCELL_X1 FILLER_0_99_241 ();
 FILLCELL_X2 FILLER_0_99_252 ();
 FILLCELL_X1 FILLER_0_99_254 ();
 FILLCELL_X4 FILLER_0_99_438 ();
 FILLCELL_X2 FILLER_0_99_481 ();
 FILLCELL_X1 FILLER_0_99_483 ();
 FILLCELL_X2 FILLER_0_99_499 ();
 FILLCELL_X1 FILLER_0_99_501 ();
 FILLCELL_X4 FILLER_0_99_551 ();
 FILLCELL_X1 FILLER_0_99_562 ();
 FILLCELL_X1 FILLER_0_99_578 ();
 FILLCELL_X16 FILLER_0_99_594 ();
 FILLCELL_X16 FILLER_0_99_623 ();
 FILLCELL_X8 FILLER_0_99_639 ();
 FILLCELL_X4 FILLER_0_99_647 ();
 FILLCELL_X1 FILLER_0_99_651 ();
 FILLCELL_X4 FILLER_0_99_656 ();
 FILLCELL_X2 FILLER_0_99_660 ();
 FILLCELL_X2 FILLER_0_99_686 ();
 FILLCELL_X2 FILLER_0_99_718 ();
 FILLCELL_X1 FILLER_0_99_720 ();
 FILLCELL_X1 FILLER_0_99_738 ();
 FILLCELL_X4 FILLER_0_99_854 ();
 FILLCELL_X2 FILLER_0_99_912 ();
 FILLCELL_X1 FILLER_0_99_914 ();
 FILLCELL_X2 FILLER_0_99_932 ();
 FILLCELL_X1 FILLER_0_99_961 ();
 FILLCELL_X1 FILLER_0_99_997 ();
 FILLCELL_X4 FILLER_0_99_1038 ();
 FILLCELL_X2 FILLER_0_99_1064 ();
 FILLCELL_X4 FILLER_0_99_1095 ();
 FILLCELL_X2 FILLER_0_99_1125 ();
 FILLCELL_X32 FILLER_0_100_1 ();
 FILLCELL_X32 FILLER_0_100_33 ();
 FILLCELL_X32 FILLER_0_100_65 ();
 FILLCELL_X32 FILLER_0_100_97 ();
 FILLCELL_X32 FILLER_0_100_129 ();
 FILLCELL_X32 FILLER_0_100_161 ();
 FILLCELL_X16 FILLER_0_100_193 ();
 FILLCELL_X1 FILLER_0_100_239 ();
 FILLCELL_X1 FILLER_0_100_261 ();
 FILLCELL_X2 FILLER_0_100_286 ();
 FILLCELL_X2 FILLER_0_100_298 ();
 FILLCELL_X1 FILLER_0_100_300 ();
 FILLCELL_X1 FILLER_0_100_328 ();
 FILLCELL_X8 FILLER_0_100_383 ();
 FILLCELL_X2 FILLER_0_100_395 ();
 FILLCELL_X1 FILLER_0_100_407 ();
 FILLCELL_X2 FILLER_0_100_415 ();
 FILLCELL_X1 FILLER_0_100_441 ();
 FILLCELL_X2 FILLER_0_100_468 ();
 FILLCELL_X1 FILLER_0_100_470 ();
 FILLCELL_X1 FILLER_0_100_490 ();
 FILLCELL_X2 FILLER_0_100_515 ();
 FILLCELL_X1 FILLER_0_100_517 ();
 FILLCELL_X2 FILLER_0_100_528 ();
 FILLCELL_X4 FILLER_0_100_569 ();
 FILLCELL_X8 FILLER_0_100_603 ();
 FILLCELL_X2 FILLER_0_100_611 ();
 FILLCELL_X1 FILLER_0_100_613 ();
 FILLCELL_X2 FILLER_0_100_619 ();
 FILLCELL_X16 FILLER_0_100_632 ();
 FILLCELL_X2 FILLER_0_100_648 ();
 FILLCELL_X1 FILLER_0_100_665 ();
 FILLCELL_X2 FILLER_0_100_721 ();
 FILLCELL_X1 FILLER_0_100_723 ();
 FILLCELL_X2 FILLER_0_100_755 ();
 FILLCELL_X2 FILLER_0_100_788 ();
 FILLCELL_X1 FILLER_0_100_817 ();
 FILLCELL_X1 FILLER_0_100_846 ();
 FILLCELL_X4 FILLER_0_100_855 ();
 FILLCELL_X2 FILLER_0_100_896 ();
 FILLCELL_X2 FILLER_0_100_928 ();
 FILLCELL_X1 FILLER_0_100_930 ();
 FILLCELL_X1 FILLER_0_100_961 ();
 FILLCELL_X1 FILLER_0_100_989 ();
 FILLCELL_X1 FILLER_0_100_1000 ();
 FILLCELL_X2 FILLER_0_100_1011 ();
 FILLCELL_X1 FILLER_0_100_1033 ();
 FILLCELL_X1 FILLER_0_100_1054 ();
 FILLCELL_X8 FILLER_0_100_1106 ();
 FILLCELL_X4 FILLER_0_100_1114 ();
 FILLCELL_X1 FILLER_0_100_1124 ();
 FILLCELL_X4 FILLER_0_101_1 ();
 FILLCELL_X2 FILLER_0_101_5 ();
 FILLCELL_X32 FILLER_0_101_32 ();
 FILLCELL_X32 FILLER_0_101_64 ();
 FILLCELL_X32 FILLER_0_101_96 ();
 FILLCELL_X32 FILLER_0_101_128 ();
 FILLCELL_X32 FILLER_0_101_160 ();
 FILLCELL_X16 FILLER_0_101_192 ();
 FILLCELL_X2 FILLER_0_101_299 ();
 FILLCELL_X1 FILLER_0_101_367 ();
 FILLCELL_X4 FILLER_0_101_385 ();
 FILLCELL_X2 FILLER_0_101_389 ();
 FILLCELL_X1 FILLER_0_101_401 ();
 FILLCELL_X4 FILLER_0_101_405 ();
 FILLCELL_X2 FILLER_0_101_409 ();
 FILLCELL_X4 FILLER_0_101_415 ();
 FILLCELL_X2 FILLER_0_101_419 ();
 FILLCELL_X1 FILLER_0_101_421 ();
 FILLCELL_X4 FILLER_0_101_432 ();
 FILLCELL_X2 FILLER_0_101_436 ();
 FILLCELL_X1 FILLER_0_101_438 ();
 FILLCELL_X1 FILLER_0_101_454 ();
 FILLCELL_X2 FILLER_0_101_498 ();
 FILLCELL_X1 FILLER_0_101_500 ();
 FILLCELL_X4 FILLER_0_101_528 ();
 FILLCELL_X2 FILLER_0_101_556 ();
 FILLCELL_X1 FILLER_0_101_558 ();
 FILLCELL_X2 FILLER_0_101_593 ();
 FILLCELL_X1 FILLER_0_101_595 ();
 FILLCELL_X2 FILLER_0_101_610 ();
 FILLCELL_X1 FILLER_0_101_612 ();
 FILLCELL_X4 FILLER_0_101_632 ();
 FILLCELL_X4 FILLER_0_101_656 ();
 FILLCELL_X1 FILLER_0_101_665 ();
 FILLCELL_X2 FILLER_0_101_686 ();
 FILLCELL_X1 FILLER_0_101_688 ();
 FILLCELL_X2 FILLER_0_101_696 ();
 FILLCELL_X1 FILLER_0_101_698 ();
 FILLCELL_X2 FILLER_0_101_734 ();
 FILLCELL_X1 FILLER_0_101_736 ();
 FILLCELL_X1 FILLER_0_101_747 ();
 FILLCELL_X1 FILLER_0_101_758 ();
 FILLCELL_X1 FILLER_0_101_769 ();
 FILLCELL_X4 FILLER_0_101_787 ();
 FILLCELL_X4 FILLER_0_101_843 ();
 FILLCELL_X2 FILLER_0_101_847 ();
 FILLCELL_X1 FILLER_0_101_849 ();
 FILLCELL_X1 FILLER_0_101_860 ();
 FILLCELL_X8 FILLER_0_101_881 ();
 FILLCELL_X4 FILLER_0_101_889 ();
 FILLCELL_X1 FILLER_0_101_907 ();
 FILLCELL_X4 FILLER_0_101_918 ();
 FILLCELL_X4 FILLER_0_101_932 ();
 FILLCELL_X1 FILLER_0_101_970 ();
 FILLCELL_X1 FILLER_0_101_981 ();
 FILLCELL_X1 FILLER_0_101_1008 ();
 FILLCELL_X2 FILLER_0_101_1026 ();
 FILLCELL_X8 FILLER_0_101_1048 ();
 FILLCELL_X4 FILLER_0_101_1056 ();
 FILLCELL_X2 FILLER_0_101_1060 ();
 FILLCELL_X32 FILLER_0_101_1087 ();
 FILLCELL_X8 FILLER_0_101_1119 ();
 FILLCELL_X8 FILLER_0_101_1130 ();
 FILLCELL_X1 FILLER_0_101_1147 ();
 FILLCELL_X32 FILLER_0_102_1 ();
 FILLCELL_X32 FILLER_0_102_33 ();
 FILLCELL_X32 FILLER_0_102_65 ();
 FILLCELL_X32 FILLER_0_102_97 ();
 FILLCELL_X32 FILLER_0_102_129 ();
 FILLCELL_X32 FILLER_0_102_161 ();
 FILLCELL_X8 FILLER_0_102_193 ();
 FILLCELL_X4 FILLER_0_102_201 ();
 FILLCELL_X1 FILLER_0_102_228 ();
 FILLCELL_X2 FILLER_0_102_253 ();
 FILLCELL_X1 FILLER_0_102_265 ();
 FILLCELL_X2 FILLER_0_102_281 ();
 FILLCELL_X1 FILLER_0_102_399 ();
 FILLCELL_X4 FILLER_0_102_407 ();
 FILLCELL_X1 FILLER_0_102_411 ();
 FILLCELL_X2 FILLER_0_102_422 ();
 FILLCELL_X2 FILLER_0_102_429 ();
 FILLCELL_X4 FILLER_0_102_441 ();
 FILLCELL_X1 FILLER_0_102_455 ();
 FILLCELL_X1 FILLER_0_102_473 ();
 FILLCELL_X2 FILLER_0_102_504 ();
 FILLCELL_X1 FILLER_0_102_506 ();
 FILLCELL_X4 FILLER_0_102_563 ();
 FILLCELL_X1 FILLER_0_102_596 ();
 FILLCELL_X4 FILLER_0_102_607 ();
 FILLCELL_X8 FILLER_0_102_632 ();
 FILLCELL_X1 FILLER_0_102_724 ();
 FILLCELL_X2 FILLER_0_102_735 ();
 FILLCELL_X1 FILLER_0_102_737 ();
 FILLCELL_X4 FILLER_0_102_798 ();
 FILLCELL_X2 FILLER_0_102_822 ();
 FILLCELL_X1 FILLER_0_102_846 ();
 FILLCELL_X1 FILLER_0_102_866 ();
 FILLCELL_X2 FILLER_0_102_884 ();
 FILLCELL_X1 FILLER_0_102_886 ();
 FILLCELL_X2 FILLER_0_102_904 ();
 FILLCELL_X4 FILLER_0_102_933 ();
 FILLCELL_X1 FILLER_0_102_944 ();
 FILLCELL_X2 FILLER_0_102_977 ();
 FILLCELL_X1 FILLER_0_102_979 ();
 FILLCELL_X2 FILLER_0_102_1011 ();
 FILLCELL_X1 FILLER_0_102_1013 ();
 FILLCELL_X1 FILLER_0_102_1024 ();
 FILLCELL_X32 FILLER_0_102_1054 ();
 FILLCELL_X32 FILLER_0_102_1086 ();
 FILLCELL_X16 FILLER_0_102_1118 ();
 FILLCELL_X8 FILLER_0_102_1134 ();
 FILLCELL_X4 FILLER_0_102_1142 ();
 FILLCELL_X2 FILLER_0_102_1146 ();
 FILLCELL_X32 FILLER_0_103_1 ();
 FILLCELL_X32 FILLER_0_103_33 ();
 FILLCELL_X32 FILLER_0_103_65 ();
 FILLCELL_X32 FILLER_0_103_97 ();
 FILLCELL_X32 FILLER_0_103_129 ();
 FILLCELL_X32 FILLER_0_103_161 ();
 FILLCELL_X8 FILLER_0_103_193 ();
 FILLCELL_X2 FILLER_0_103_201 ();
 FILLCELL_X1 FILLER_0_103_307 ();
 FILLCELL_X2 FILLER_0_103_365 ();
 FILLCELL_X4 FILLER_0_103_388 ();
 FILLCELL_X4 FILLER_0_103_433 ();
 FILLCELL_X2 FILLER_0_103_551 ();
 FILLCELL_X1 FILLER_0_103_604 ();
 FILLCELL_X8 FILLER_0_103_615 ();
 FILLCELL_X4 FILLER_0_103_623 ();
 FILLCELL_X2 FILLER_0_103_637 ();
 FILLCELL_X1 FILLER_0_103_639 ();
 FILLCELL_X1 FILLER_0_103_673 ();
 FILLCELL_X1 FILLER_0_103_691 ();
 FILLCELL_X1 FILLER_0_103_716 ();
 FILLCELL_X1 FILLER_0_103_734 ();
 FILLCELL_X1 FILLER_0_103_745 ();
 FILLCELL_X2 FILLER_0_103_777 ();
 FILLCELL_X1 FILLER_0_103_779 ();
 FILLCELL_X4 FILLER_0_103_815 ();
 FILLCELL_X2 FILLER_0_103_819 ();
 FILLCELL_X1 FILLER_0_103_821 ();
 FILLCELL_X4 FILLER_0_103_827 ();
 FILLCELL_X2 FILLER_0_103_855 ();
 FILLCELL_X1 FILLER_0_103_857 ();
 FILLCELL_X2 FILLER_0_103_867 ();
 FILLCELL_X4 FILLER_0_103_893 ();
 FILLCELL_X1 FILLER_0_103_902 ();
 FILLCELL_X1 FILLER_0_103_927 ();
 FILLCELL_X1 FILLER_0_103_942 ();
 FILLCELL_X1 FILLER_0_103_957 ();
 FILLCELL_X1 FILLER_0_103_968 ();
 FILLCELL_X1 FILLER_0_103_979 ();
 FILLCELL_X1 FILLER_0_103_1002 ();
 FILLCELL_X4 FILLER_0_103_1020 ();
 FILLCELL_X2 FILLER_0_103_1040 ();
 FILLCELL_X1 FILLER_0_103_1042 ();
 FILLCELL_X32 FILLER_0_103_1063 ();
 FILLCELL_X32 FILLER_0_103_1095 ();
 FILLCELL_X16 FILLER_0_103_1127 ();
 FILLCELL_X4 FILLER_0_103_1143 ();
 FILLCELL_X1 FILLER_0_103_1147 ();
 FILLCELL_X32 FILLER_0_104_1 ();
 FILLCELL_X32 FILLER_0_104_33 ();
 FILLCELL_X32 FILLER_0_104_65 ();
 FILLCELL_X32 FILLER_0_104_97 ();
 FILLCELL_X32 FILLER_0_104_129 ();
 FILLCELL_X32 FILLER_0_104_161 ();
 FILLCELL_X8 FILLER_0_104_193 ();
 FILLCELL_X4 FILLER_0_104_201 ();
 FILLCELL_X2 FILLER_0_104_205 ();
 FILLCELL_X1 FILLER_0_104_207 ();
 FILLCELL_X1 FILLER_0_104_244 ();
 FILLCELL_X2 FILLER_0_104_262 ();
 FILLCELL_X2 FILLER_0_104_295 ();
 FILLCELL_X1 FILLER_0_104_297 ();
 FILLCELL_X2 FILLER_0_104_308 ();
 FILLCELL_X1 FILLER_0_104_337 ();
 FILLCELL_X1 FILLER_0_104_348 ();
 FILLCELL_X1 FILLER_0_104_366 ();
 FILLCELL_X4 FILLER_0_104_415 ();
 FILLCELL_X2 FILLER_0_104_419 ();
 FILLCELL_X4 FILLER_0_104_474 ();
 FILLCELL_X2 FILLER_0_104_502 ();
 FILLCELL_X1 FILLER_0_104_504 ();
 FILLCELL_X2 FILLER_0_104_532 ();
 FILLCELL_X2 FILLER_0_104_551 ();
 FILLCELL_X1 FILLER_0_104_553 ();
 FILLCELL_X2 FILLER_0_104_564 ();
 FILLCELL_X1 FILLER_0_104_630 ();
 FILLCELL_X16 FILLER_0_104_632 ();
 FILLCELL_X4 FILLER_0_104_648 ();
 FILLCELL_X2 FILLER_0_104_659 ();
 FILLCELL_X1 FILLER_0_104_676 ();
 FILLCELL_X1 FILLER_0_104_703 ();
 FILLCELL_X1 FILLER_0_104_725 ();
 FILLCELL_X2 FILLER_0_104_740 ();
 FILLCELL_X1 FILLER_0_104_752 ();
 FILLCELL_X1 FILLER_0_104_763 ();
 FILLCELL_X4 FILLER_0_104_795 ();
 FILLCELL_X16 FILLER_0_104_814 ();
 FILLCELL_X4 FILLER_0_104_830 ();
 FILLCELL_X2 FILLER_0_104_834 ();
 FILLCELL_X4 FILLER_0_104_850 ();
 FILLCELL_X1 FILLER_0_104_854 ();
 FILLCELL_X8 FILLER_0_104_865 ();
 FILLCELL_X1 FILLER_0_104_873 ();
 FILLCELL_X4 FILLER_0_104_884 ();
 FILLCELL_X1 FILLER_0_104_898 ();
 FILLCELL_X1 FILLER_0_104_909 ();
 FILLCELL_X2 FILLER_0_104_924 ();
 FILLCELL_X1 FILLER_0_104_926 ();
 FILLCELL_X4 FILLER_0_104_941 ();
 FILLCELL_X4 FILLER_0_104_977 ();
 FILLCELL_X4 FILLER_0_104_1010 ();
 FILLCELL_X32 FILLER_0_104_1054 ();
 FILLCELL_X32 FILLER_0_104_1086 ();
 FILLCELL_X16 FILLER_0_104_1118 ();
 FILLCELL_X8 FILLER_0_104_1134 ();
 FILLCELL_X4 FILLER_0_104_1142 ();
 FILLCELL_X2 FILLER_0_104_1146 ();
 FILLCELL_X32 FILLER_0_105_1 ();
 FILLCELL_X32 FILLER_0_105_33 ();
 FILLCELL_X32 FILLER_0_105_65 ();
 FILLCELL_X32 FILLER_0_105_97 ();
 FILLCELL_X32 FILLER_0_105_129 ();
 FILLCELL_X32 FILLER_0_105_161 ();
 FILLCELL_X16 FILLER_0_105_193 ();
 FILLCELL_X2 FILLER_0_105_209 ();
 FILLCELL_X1 FILLER_0_105_211 ();
 FILLCELL_X4 FILLER_0_105_230 ();
 FILLCELL_X4 FILLER_0_105_273 ();
 FILLCELL_X1 FILLER_0_105_331 ();
 FILLCELL_X2 FILLER_0_105_342 ();
 FILLCELL_X1 FILLER_0_105_354 ();
 FILLCELL_X16 FILLER_0_105_387 ();
 FILLCELL_X8 FILLER_0_105_412 ();
 FILLCELL_X4 FILLER_0_105_420 ();
 FILLCELL_X1 FILLER_0_105_434 ();
 FILLCELL_X1 FILLER_0_105_445 ();
 FILLCELL_X1 FILLER_0_105_456 ();
 FILLCELL_X2 FILLER_0_105_472 ();
 FILLCELL_X2 FILLER_0_105_501 ();
 FILLCELL_X1 FILLER_0_105_503 ();
 FILLCELL_X2 FILLER_0_105_524 ();
 FILLCELL_X1 FILLER_0_105_526 ();
 FILLCELL_X2 FILLER_0_105_537 ();
 FILLCELL_X2 FILLER_0_105_556 ();
 FILLCELL_X2 FILLER_0_105_598 ();
 FILLCELL_X1 FILLER_0_105_600 ();
 FILLCELL_X16 FILLER_0_105_616 ();
 FILLCELL_X4 FILLER_0_105_632 ();
 FILLCELL_X2 FILLER_0_105_636 ();
 FILLCELL_X1 FILLER_0_105_638 ();
 FILLCELL_X2 FILLER_0_105_653 ();
 FILLCELL_X2 FILLER_0_105_674 ();
 FILLCELL_X2 FILLER_0_105_686 ();
 FILLCELL_X1 FILLER_0_105_688 ();
 FILLCELL_X2 FILLER_0_105_758 ();
 FILLCELL_X1 FILLER_0_105_760 ();
 FILLCELL_X4 FILLER_0_105_770 ();
 FILLCELL_X4 FILLER_0_105_783 ();
 FILLCELL_X1 FILLER_0_105_852 ();
 FILLCELL_X1 FILLER_0_105_858 ();
 FILLCELL_X2 FILLER_0_105_868 ();
 FILLCELL_X1 FILLER_0_105_884 ();
 FILLCELL_X1 FILLER_0_105_900 ();
 FILLCELL_X2 FILLER_0_105_911 ();
 FILLCELL_X1 FILLER_0_105_933 ();
 FILLCELL_X2 FILLER_0_105_958 ();
 FILLCELL_X1 FILLER_0_105_975 ();
 FILLCELL_X2 FILLER_0_105_993 ();
 FILLCELL_X4 FILLER_0_105_1005 ();
 FILLCELL_X4 FILLER_0_105_1049 ();
 FILLCELL_X1 FILLER_0_105_1053 ();
 FILLCELL_X32 FILLER_0_105_1064 ();
 FILLCELL_X32 FILLER_0_105_1096 ();
 FILLCELL_X16 FILLER_0_105_1128 ();
 FILLCELL_X4 FILLER_0_105_1144 ();
 FILLCELL_X32 FILLER_0_106_1 ();
 FILLCELL_X32 FILLER_0_106_33 ();
 FILLCELL_X32 FILLER_0_106_65 ();
 FILLCELL_X32 FILLER_0_106_97 ();
 FILLCELL_X32 FILLER_0_106_129 ();
 FILLCELL_X32 FILLER_0_106_161 ();
 FILLCELL_X16 FILLER_0_106_193 ();
 FILLCELL_X4 FILLER_0_106_209 ();
 FILLCELL_X1 FILLER_0_106_289 ();
 FILLCELL_X1 FILLER_0_106_353 ();
 FILLCELL_X16 FILLER_0_106_418 ();
 FILLCELL_X4 FILLER_0_106_434 ();
 FILLCELL_X2 FILLER_0_106_438 ();
 FILLCELL_X1 FILLER_0_106_440 ();
 FILLCELL_X4 FILLER_0_106_451 ();
 FILLCELL_X2 FILLER_0_106_465 ();
 FILLCELL_X1 FILLER_0_106_467 ();
 FILLCELL_X1 FILLER_0_106_475 ();
 FILLCELL_X2 FILLER_0_106_514 ();
 FILLCELL_X2 FILLER_0_106_533 ();
 FILLCELL_X2 FILLER_0_106_549 ();
 FILLCELL_X1 FILLER_0_106_590 ();
 FILLCELL_X1 FILLER_0_106_601 ();
 FILLCELL_X4 FILLER_0_106_626 ();
 FILLCELL_X1 FILLER_0_106_630 ();
 FILLCELL_X8 FILLER_0_106_632 ();
 FILLCELL_X2 FILLER_0_106_640 ();
 FILLCELL_X1 FILLER_0_106_642 ();
 FILLCELL_X2 FILLER_0_106_683 ();
 FILLCELL_X2 FILLER_0_106_692 ();
 FILLCELL_X1 FILLER_0_106_694 ();
 FILLCELL_X1 FILLER_0_106_710 ();
 FILLCELL_X2 FILLER_0_106_721 ();
 FILLCELL_X1 FILLER_0_106_723 ();
 FILLCELL_X1 FILLER_0_106_776 ();
 FILLCELL_X1 FILLER_0_106_804 ();
 FILLCELL_X2 FILLER_0_106_820 ();
 FILLCELL_X2 FILLER_0_106_832 ();
 FILLCELL_X1 FILLER_0_106_834 ();
 FILLCELL_X1 FILLER_0_106_845 ();
 FILLCELL_X1 FILLER_0_106_914 ();
 FILLCELL_X2 FILLER_0_106_940 ();
 FILLCELL_X1 FILLER_0_106_978 ();
 FILLCELL_X2 FILLER_0_106_1028 ();
 FILLCELL_X32 FILLER_0_106_1050 ();
 FILLCELL_X32 FILLER_0_106_1082 ();
 FILLCELL_X32 FILLER_0_106_1114 ();
 FILLCELL_X2 FILLER_0_106_1146 ();
 FILLCELL_X32 FILLER_0_107_1 ();
 FILLCELL_X32 FILLER_0_107_33 ();
 FILLCELL_X32 FILLER_0_107_65 ();
 FILLCELL_X32 FILLER_0_107_97 ();
 FILLCELL_X32 FILLER_0_107_129 ();
 FILLCELL_X32 FILLER_0_107_161 ();
 FILLCELL_X8 FILLER_0_107_193 ();
 FILLCELL_X4 FILLER_0_107_201 ();
 FILLCELL_X1 FILLER_0_107_205 ();
 FILLCELL_X1 FILLER_0_107_234 ();
 FILLCELL_X1 FILLER_0_107_245 ();
 FILLCELL_X1 FILLER_0_107_255 ();
 FILLCELL_X1 FILLER_0_107_286 ();
 FILLCELL_X2 FILLER_0_107_319 ();
 FILLCELL_X1 FILLER_0_107_328 ();
 FILLCELL_X1 FILLER_0_107_354 ();
 FILLCELL_X1 FILLER_0_107_370 ();
 FILLCELL_X8 FILLER_0_107_392 ();
 FILLCELL_X2 FILLER_0_107_400 ();
 FILLCELL_X1 FILLER_0_107_402 ();
 FILLCELL_X2 FILLER_0_107_412 ();
 FILLCELL_X16 FILLER_0_107_429 ();
 FILLCELL_X4 FILLER_0_107_445 ();
 FILLCELL_X1 FILLER_0_107_449 ();
 FILLCELL_X4 FILLER_0_107_470 ();
 FILLCELL_X2 FILLER_0_107_499 ();
 FILLCELL_X2 FILLER_0_107_544 ();
 FILLCELL_X1 FILLER_0_107_556 ();
 FILLCELL_X1 FILLER_0_107_567 ();
 FILLCELL_X1 FILLER_0_107_573 ();
 FILLCELL_X1 FILLER_0_107_584 ();
 FILLCELL_X2 FILLER_0_107_595 ();
 FILLCELL_X1 FILLER_0_107_607 ();
 FILLCELL_X2 FILLER_0_107_613 ();
 FILLCELL_X2 FILLER_0_107_625 ();
 FILLCELL_X4 FILLER_0_107_637 ();
 FILLCELL_X4 FILLER_0_107_723 ();
 FILLCELL_X1 FILLER_0_107_742 ();
 FILLCELL_X2 FILLER_0_107_767 ();
 FILLCELL_X1 FILLER_0_107_779 ();
 FILLCELL_X4 FILLER_0_107_790 ();
 FILLCELL_X1 FILLER_0_107_809 ();
 FILLCELL_X2 FILLER_0_107_815 ();
 FILLCELL_X1 FILLER_0_107_817 ();
 FILLCELL_X8 FILLER_0_107_828 ();
 FILLCELL_X4 FILLER_0_107_836 ();
 FILLCELL_X2 FILLER_0_107_840 ();
 FILLCELL_X1 FILLER_0_107_842 ();
 FILLCELL_X8 FILLER_0_107_853 ();
 FILLCELL_X2 FILLER_0_107_876 ();
 FILLCELL_X1 FILLER_0_107_878 ();
 FILLCELL_X4 FILLER_0_107_928 ();
 FILLCELL_X2 FILLER_0_107_949 ();
 FILLCELL_X1 FILLER_0_107_951 ();
 FILLCELL_X2 FILLER_0_107_962 ();
 FILLCELL_X4 FILLER_0_107_971 ();
 FILLCELL_X2 FILLER_0_107_992 ();
 FILLCELL_X1 FILLER_0_107_994 ();
 FILLCELL_X2 FILLER_0_107_1040 ();
 FILLCELL_X1 FILLER_0_107_1042 ();
 FILLCELL_X32 FILLER_0_107_1063 ();
 FILLCELL_X32 FILLER_0_107_1095 ();
 FILLCELL_X16 FILLER_0_107_1127 ();
 FILLCELL_X4 FILLER_0_107_1143 ();
 FILLCELL_X1 FILLER_0_107_1147 ();
 FILLCELL_X32 FILLER_0_108_1 ();
 FILLCELL_X32 FILLER_0_108_33 ();
 FILLCELL_X32 FILLER_0_108_65 ();
 FILLCELL_X32 FILLER_0_108_97 ();
 FILLCELL_X32 FILLER_0_108_129 ();
 FILLCELL_X32 FILLER_0_108_161 ();
 FILLCELL_X32 FILLER_0_108_193 ();
 FILLCELL_X2 FILLER_0_108_225 ();
 FILLCELL_X1 FILLER_0_108_227 ();
 FILLCELL_X1 FILLER_0_108_243 ();
 FILLCELL_X1 FILLER_0_108_254 ();
 FILLCELL_X1 FILLER_0_108_264 ();
 FILLCELL_X4 FILLER_0_108_342 ();
 FILLCELL_X1 FILLER_0_108_355 ();
 FILLCELL_X2 FILLER_0_108_383 ();
 FILLCELL_X1 FILLER_0_108_385 ();
 FILLCELL_X4 FILLER_0_108_396 ();
 FILLCELL_X2 FILLER_0_108_400 ();
 FILLCELL_X1 FILLER_0_108_439 ();
 FILLCELL_X4 FILLER_0_108_464 ();
 FILLCELL_X2 FILLER_0_108_475 ();
 FILLCELL_X1 FILLER_0_108_477 ();
 FILLCELL_X2 FILLER_0_108_503 ();
 FILLCELL_X1 FILLER_0_108_505 ();
 FILLCELL_X8 FILLER_0_108_594 ();
 FILLCELL_X4 FILLER_0_108_602 ();
 FILLCELL_X1 FILLER_0_108_606 ();
 FILLCELL_X4 FILLER_0_108_627 ();
 FILLCELL_X8 FILLER_0_108_632 ();
 FILLCELL_X4 FILLER_0_108_640 ();
 FILLCELL_X1 FILLER_0_108_644 ();
 FILLCELL_X2 FILLER_0_108_655 ();
 FILLCELL_X1 FILLER_0_108_657 ();
 FILLCELL_X4 FILLER_0_108_668 ();
 FILLCELL_X2 FILLER_0_108_672 ();
 FILLCELL_X2 FILLER_0_108_716 ();
 FILLCELL_X1 FILLER_0_108_735 ();
 FILLCELL_X4 FILLER_0_108_750 ();
 FILLCELL_X4 FILLER_0_108_771 ();
 FILLCELL_X2 FILLER_0_108_792 ();
 FILLCELL_X1 FILLER_0_108_794 ();
 FILLCELL_X2 FILLER_0_108_805 ();
 FILLCELL_X1 FILLER_0_108_807 ();
 FILLCELL_X16 FILLER_0_108_818 ();
 FILLCELL_X2 FILLER_0_108_834 ();
 FILLCELL_X2 FILLER_0_108_853 ();
 FILLCELL_X1 FILLER_0_108_855 ();
 FILLCELL_X2 FILLER_0_108_918 ();
 FILLCELL_X1 FILLER_0_108_959 ();
 FILLCELL_X1 FILLER_0_108_970 ();
 FILLCELL_X2 FILLER_0_108_985 ();
 FILLCELL_X4 FILLER_0_108_1022 ();
 FILLCELL_X1 FILLER_0_108_1026 ();
 FILLCELL_X2 FILLER_0_108_1037 ();
 FILLCELL_X32 FILLER_0_108_1064 ();
 FILLCELL_X32 FILLER_0_108_1096 ();
 FILLCELL_X16 FILLER_0_108_1128 ();
 FILLCELL_X4 FILLER_0_108_1144 ();
 FILLCELL_X32 FILLER_0_109_1 ();
 FILLCELL_X32 FILLER_0_109_33 ();
 FILLCELL_X32 FILLER_0_109_65 ();
 FILLCELL_X32 FILLER_0_109_97 ();
 FILLCELL_X32 FILLER_0_109_129 ();
 FILLCELL_X32 FILLER_0_109_161 ();
 FILLCELL_X16 FILLER_0_109_193 ();
 FILLCELL_X8 FILLER_0_109_209 ();
 FILLCELL_X4 FILLER_0_109_217 ();
 FILLCELL_X2 FILLER_0_109_221 ();
 FILLCELL_X2 FILLER_0_109_235 ();
 FILLCELL_X1 FILLER_0_109_247 ();
 FILLCELL_X1 FILLER_0_109_273 ();
 FILLCELL_X1 FILLER_0_109_301 ();
 FILLCELL_X2 FILLER_0_109_375 ();
 FILLCELL_X2 FILLER_0_109_397 ();
 FILLCELL_X1 FILLER_0_109_414 ();
 FILLCELL_X1 FILLER_0_109_425 ();
 FILLCELL_X1 FILLER_0_109_431 ();
 FILLCELL_X4 FILLER_0_109_451 ();
 FILLCELL_X1 FILLER_0_109_455 ();
 FILLCELL_X2 FILLER_0_109_483 ();
 FILLCELL_X1 FILLER_0_109_495 ();
 FILLCELL_X1 FILLER_0_109_505 ();
 FILLCELL_X1 FILLER_0_109_520 ();
 FILLCELL_X1 FILLER_0_109_538 ();
 FILLCELL_X2 FILLER_0_109_578 ();
 FILLCELL_X16 FILLER_0_109_590 ();
 FILLCELL_X4 FILLER_0_109_606 ();
 FILLCELL_X1 FILLER_0_109_610 ();
 FILLCELL_X16 FILLER_0_109_621 ();
 FILLCELL_X8 FILLER_0_109_637 ();
 FILLCELL_X4 FILLER_0_109_645 ();
 FILLCELL_X2 FILLER_0_109_649 ();
 FILLCELL_X1 FILLER_0_109_651 ();
 FILLCELL_X8 FILLER_0_109_671 ();
 FILLCELL_X2 FILLER_0_109_679 ();
 FILLCELL_X2 FILLER_0_109_691 ();
 FILLCELL_X1 FILLER_0_109_693 ();
 FILLCELL_X2 FILLER_0_109_709 ();
 FILLCELL_X1 FILLER_0_109_721 ();
 FILLCELL_X1 FILLER_0_109_746 ();
 FILLCELL_X1 FILLER_0_109_762 ();
 FILLCELL_X1 FILLER_0_109_770 ();
 FILLCELL_X2 FILLER_0_109_803 ();
 FILLCELL_X1 FILLER_0_109_805 ();
 FILLCELL_X8 FILLER_0_109_821 ();
 FILLCELL_X2 FILLER_0_109_829 ();
 FILLCELL_X4 FILLER_0_109_841 ();
 FILLCELL_X2 FILLER_0_109_845 ();
 FILLCELL_X1 FILLER_0_109_847 ();
 FILLCELL_X4 FILLER_0_109_853 ();
 FILLCELL_X1 FILLER_0_109_857 ();
 FILLCELL_X4 FILLER_0_109_863 ();
 FILLCELL_X2 FILLER_0_109_867 ();
 FILLCELL_X1 FILLER_0_109_869 ();
 FILLCELL_X1 FILLER_0_109_909 ();
 FILLCELL_X1 FILLER_0_109_939 ();
 FILLCELL_X4 FILLER_0_109_969 ();
 FILLCELL_X1 FILLER_0_109_998 ();
 FILLCELL_X2 FILLER_0_109_1019 ();
 FILLCELL_X4 FILLER_0_109_1031 ();
 FILLCELL_X32 FILLER_0_109_1054 ();
 FILLCELL_X32 FILLER_0_109_1086 ();
 FILLCELL_X16 FILLER_0_109_1118 ();
 FILLCELL_X8 FILLER_0_109_1134 ();
 FILLCELL_X4 FILLER_0_109_1142 ();
 FILLCELL_X2 FILLER_0_109_1146 ();
 FILLCELL_X32 FILLER_0_110_1 ();
 FILLCELL_X32 FILLER_0_110_33 ();
 FILLCELL_X32 FILLER_0_110_65 ();
 FILLCELL_X32 FILLER_0_110_97 ();
 FILLCELL_X32 FILLER_0_110_129 ();
 FILLCELL_X32 FILLER_0_110_161 ();
 FILLCELL_X16 FILLER_0_110_193 ();
 FILLCELL_X1 FILLER_0_110_209 ();
 FILLCELL_X1 FILLER_0_110_219 ();
 FILLCELL_X2 FILLER_0_110_238 ();
 FILLCELL_X2 FILLER_0_110_250 ();
 FILLCELL_X2 FILLER_0_110_267 ();
 FILLCELL_X1 FILLER_0_110_279 ();
 FILLCELL_X2 FILLER_0_110_296 ();
 FILLCELL_X1 FILLER_0_110_298 ();
 FILLCELL_X1 FILLER_0_110_306 ();
 FILLCELL_X2 FILLER_0_110_324 ();
 FILLCELL_X1 FILLER_0_110_326 ();
 FILLCELL_X2 FILLER_0_110_337 ();
 FILLCELL_X1 FILLER_0_110_339 ();
 FILLCELL_X2 FILLER_0_110_350 ();
 FILLCELL_X2 FILLER_0_110_367 ();
 FILLCELL_X2 FILLER_0_110_374 ();
 FILLCELL_X1 FILLER_0_110_376 ();
 FILLCELL_X8 FILLER_0_110_387 ();
 FILLCELL_X4 FILLER_0_110_395 ();
 FILLCELL_X1 FILLER_0_110_399 ();
 FILLCELL_X2 FILLER_0_110_410 ();
 FILLCELL_X2 FILLER_0_110_421 ();
 FILLCELL_X1 FILLER_0_110_423 ();
 FILLCELL_X8 FILLER_0_110_434 ();
 FILLCELL_X4 FILLER_0_110_442 ();
 FILLCELL_X2 FILLER_0_110_446 ();
 FILLCELL_X1 FILLER_0_110_458 ();
 FILLCELL_X2 FILLER_0_110_484 ();
 FILLCELL_X2 FILLER_0_110_515 ();
 FILLCELL_X1 FILLER_0_110_517 ();
 FILLCELL_X2 FILLER_0_110_538 ();
 FILLCELL_X1 FILLER_0_110_540 ();
 FILLCELL_X1 FILLER_0_110_586 ();
 FILLCELL_X4 FILLER_0_110_592 ();
 FILLCELL_X1 FILLER_0_110_606 ();
 FILLCELL_X2 FILLER_0_110_617 ();
 FILLCELL_X2 FILLER_0_110_629 ();
 FILLCELL_X8 FILLER_0_110_632 ();
 FILLCELL_X1 FILLER_0_110_640 ();
 FILLCELL_X2 FILLER_0_110_666 ();
 FILLCELL_X8 FILLER_0_110_678 ();
 FILLCELL_X2 FILLER_0_110_686 ();
 FILLCELL_X1 FILLER_0_110_688 ();
 FILLCELL_X4 FILLER_0_110_696 ();
 FILLCELL_X1 FILLER_0_110_700 ();
 FILLCELL_X2 FILLER_0_110_716 ();
 FILLCELL_X2 FILLER_0_110_742 ();
 FILLCELL_X4 FILLER_0_110_786 ();
 FILLCELL_X2 FILLER_0_110_790 ();
 FILLCELL_X1 FILLER_0_110_792 ();
 FILLCELL_X2 FILLER_0_110_803 ();
 FILLCELL_X16 FILLER_0_110_815 ();
 FILLCELL_X4 FILLER_0_110_836 ();
 FILLCELL_X2 FILLER_0_110_855 ();
 FILLCELL_X4 FILLER_0_110_867 ();
 FILLCELL_X1 FILLER_0_110_871 ();
 FILLCELL_X4 FILLER_0_110_882 ();
 FILLCELL_X2 FILLER_0_110_944 ();
 FILLCELL_X1 FILLER_0_110_946 ();
 FILLCELL_X2 FILLER_0_110_966 ();
 FILLCELL_X1 FILLER_0_110_968 ();
 FILLCELL_X2 FILLER_0_110_1004 ();
 FILLCELL_X32 FILLER_0_110_1045 ();
 FILLCELL_X32 FILLER_0_110_1077 ();
 FILLCELL_X32 FILLER_0_110_1109 ();
 FILLCELL_X4 FILLER_0_110_1141 ();
 FILLCELL_X2 FILLER_0_110_1145 ();
 FILLCELL_X1 FILLER_0_110_1147 ();
 FILLCELL_X32 FILLER_0_111_1 ();
 FILLCELL_X32 FILLER_0_111_33 ();
 FILLCELL_X32 FILLER_0_111_65 ();
 FILLCELL_X32 FILLER_0_111_97 ();
 FILLCELL_X32 FILLER_0_111_129 ();
 FILLCELL_X32 FILLER_0_111_161 ();
 FILLCELL_X8 FILLER_0_111_193 ();
 FILLCELL_X4 FILLER_0_111_201 ();
 FILLCELL_X1 FILLER_0_111_215 ();
 FILLCELL_X1 FILLER_0_111_235 ();
 FILLCELL_X4 FILLER_0_111_245 ();
 FILLCELL_X2 FILLER_0_111_268 ();
 FILLCELL_X4 FILLER_0_111_280 ();
 FILLCELL_X2 FILLER_0_111_291 ();
 FILLCELL_X1 FILLER_0_111_303 ();
 FILLCELL_X2 FILLER_0_111_309 ();
 FILLCELL_X2 FILLER_0_111_333 ();
 FILLCELL_X16 FILLER_0_111_355 ();
 FILLCELL_X8 FILLER_0_111_376 ();
 FILLCELL_X4 FILLER_0_111_384 ();
 FILLCELL_X2 FILLER_0_111_388 ();
 FILLCELL_X8 FILLER_0_111_399 ();
 FILLCELL_X1 FILLER_0_111_407 ();
 FILLCELL_X4 FILLER_0_111_433 ();
 FILLCELL_X2 FILLER_0_111_437 ();
 FILLCELL_X1 FILLER_0_111_439 ();
 FILLCELL_X8 FILLER_0_111_450 ();
 FILLCELL_X2 FILLER_0_111_458 ();
 FILLCELL_X1 FILLER_0_111_469 ();
 FILLCELL_X2 FILLER_0_111_499 ();
 FILLCELL_X1 FILLER_0_111_501 ();
 FILLCELL_X2 FILLER_0_111_512 ();
 FILLCELL_X1 FILLER_0_111_519 ();
 FILLCELL_X4 FILLER_0_111_530 ();
 FILLCELL_X4 FILLER_0_111_544 ();
 FILLCELL_X2 FILLER_0_111_597 ();
 FILLCELL_X1 FILLER_0_111_639 ();
 FILLCELL_X8 FILLER_0_111_650 ();
 FILLCELL_X4 FILLER_0_111_663 ();
 FILLCELL_X2 FILLER_0_111_667 ();
 FILLCELL_X1 FILLER_0_111_669 ();
 FILLCELL_X4 FILLER_0_111_675 ();
 FILLCELL_X1 FILLER_0_111_679 ();
 FILLCELL_X4 FILLER_0_111_700 ();
 FILLCELL_X2 FILLER_0_111_714 ();
 FILLCELL_X2 FILLER_0_111_721 ();
 FILLCELL_X1 FILLER_0_111_723 ();
 FILLCELL_X2 FILLER_0_111_729 ();
 FILLCELL_X2 FILLER_0_111_751 ();
 FILLCELL_X1 FILLER_0_111_777 ();
 FILLCELL_X2 FILLER_0_111_798 ();
 FILLCELL_X16 FILLER_0_111_810 ();
 FILLCELL_X2 FILLER_0_111_836 ();
 FILLCELL_X1 FILLER_0_111_868 ();
 FILLCELL_X2 FILLER_0_111_874 ();
 FILLCELL_X2 FILLER_0_111_923 ();
 FILLCELL_X1 FILLER_0_111_925 ();
 FILLCELL_X2 FILLER_0_111_936 ();
 FILLCELL_X1 FILLER_0_111_938 ();
 FILLCELL_X2 FILLER_0_111_954 ();
 FILLCELL_X2 FILLER_0_111_991 ();
 FILLCELL_X2 FILLER_0_111_1003 ();
 FILLCELL_X1 FILLER_0_111_1005 ();
 FILLCELL_X1 FILLER_0_111_1036 ();
 FILLCELL_X32 FILLER_0_111_1047 ();
 FILLCELL_X32 FILLER_0_111_1079 ();
 FILLCELL_X32 FILLER_0_111_1111 ();
 FILLCELL_X4 FILLER_0_111_1143 ();
 FILLCELL_X1 FILLER_0_111_1147 ();
 FILLCELL_X32 FILLER_0_112_1 ();
 FILLCELL_X32 FILLER_0_112_33 ();
 FILLCELL_X32 FILLER_0_112_65 ();
 FILLCELL_X32 FILLER_0_112_97 ();
 FILLCELL_X32 FILLER_0_112_129 ();
 FILLCELL_X32 FILLER_0_112_161 ();
 FILLCELL_X16 FILLER_0_112_193 ();
 FILLCELL_X4 FILLER_0_112_209 ();
 FILLCELL_X1 FILLER_0_112_213 ();
 FILLCELL_X2 FILLER_0_112_224 ();
 FILLCELL_X2 FILLER_0_112_235 ();
 FILLCELL_X1 FILLER_0_112_237 ();
 FILLCELL_X1 FILLER_0_112_248 ();
 FILLCELL_X2 FILLER_0_112_267 ();
 FILLCELL_X1 FILLER_0_112_269 ();
 FILLCELL_X4 FILLER_0_112_289 ();
 FILLCELL_X1 FILLER_0_112_303 ();
 FILLCELL_X1 FILLER_0_112_314 ();
 FILLCELL_X4 FILLER_0_112_344 ();
 FILLCELL_X1 FILLER_0_112_348 ();
 FILLCELL_X1 FILLER_0_112_374 ();
 FILLCELL_X1 FILLER_0_112_380 ();
 FILLCELL_X1 FILLER_0_112_391 ();
 FILLCELL_X1 FILLER_0_112_397 ();
 FILLCELL_X8 FILLER_0_112_408 ();
 FILLCELL_X2 FILLER_0_112_416 ();
 FILLCELL_X1 FILLER_0_112_418 ();
 FILLCELL_X8 FILLER_0_112_429 ();
 FILLCELL_X2 FILLER_0_112_437 ();
 FILLCELL_X1 FILLER_0_112_439 ();
 FILLCELL_X8 FILLER_0_112_450 ();
 FILLCELL_X2 FILLER_0_112_458 ();
 FILLCELL_X1 FILLER_0_112_460 ();
 FILLCELL_X2 FILLER_0_112_471 ();
 FILLCELL_X1 FILLER_0_112_473 ();
 FILLCELL_X1 FILLER_0_112_484 ();
 FILLCELL_X1 FILLER_0_112_515 ();
 FILLCELL_X1 FILLER_0_112_521 ();
 FILLCELL_X2 FILLER_0_112_532 ();
 FILLCELL_X1 FILLER_0_112_534 ();
 FILLCELL_X1 FILLER_0_112_540 ();
 FILLCELL_X4 FILLER_0_112_580 ();
 FILLCELL_X1 FILLER_0_112_603 ();
 FILLCELL_X2 FILLER_0_112_609 ();
 FILLCELL_X1 FILLER_0_112_611 ();
 FILLCELL_X16 FILLER_0_112_632 ();
 FILLCELL_X2 FILLER_0_112_648 ();
 FILLCELL_X2 FILLER_0_112_670 ();
 FILLCELL_X4 FILLER_0_112_682 ();
 FILLCELL_X1 FILLER_0_112_686 ();
 FILLCELL_X4 FILLER_0_112_706 ();
 FILLCELL_X2 FILLER_0_112_710 ();
 FILLCELL_X4 FILLER_0_112_727 ();
 FILLCELL_X2 FILLER_0_112_746 ();
 FILLCELL_X1 FILLER_0_112_748 ();
 FILLCELL_X1 FILLER_0_112_754 ();
 FILLCELL_X4 FILLER_0_112_770 ();
 FILLCELL_X2 FILLER_0_112_774 ();
 FILLCELL_X8 FILLER_0_112_816 ();
 FILLCELL_X2 FILLER_0_112_843 ();
 FILLCELL_X1 FILLER_0_112_854 ();
 FILLCELL_X2 FILLER_0_112_880 ();
 FILLCELL_X4 FILLER_0_112_897 ();
 FILLCELL_X4 FILLER_0_112_916 ();
 FILLCELL_X4 FILLER_0_112_940 ();
 FILLCELL_X2 FILLER_0_112_954 ();
 FILLCELL_X1 FILLER_0_112_956 ();
 FILLCELL_X2 FILLER_0_112_991 ();
 FILLCELL_X1 FILLER_0_112_993 ();
 FILLCELL_X4 FILLER_0_112_1018 ();
 FILLCELL_X32 FILLER_0_112_1042 ();
 FILLCELL_X32 FILLER_0_112_1074 ();
 FILLCELL_X32 FILLER_0_112_1106 ();
 FILLCELL_X8 FILLER_0_112_1138 ();
 FILLCELL_X2 FILLER_0_112_1146 ();
 FILLCELL_X32 FILLER_0_113_1 ();
 FILLCELL_X32 FILLER_0_113_33 ();
 FILLCELL_X32 FILLER_0_113_65 ();
 FILLCELL_X32 FILLER_0_113_97 ();
 FILLCELL_X32 FILLER_0_113_129 ();
 FILLCELL_X32 FILLER_0_113_161 ();
 FILLCELL_X16 FILLER_0_113_193 ();
 FILLCELL_X1 FILLER_0_113_209 ();
 FILLCELL_X2 FILLER_0_113_230 ();
 FILLCELL_X1 FILLER_0_113_232 ();
 FILLCELL_X2 FILLER_0_113_271 ();
 FILLCELL_X2 FILLER_0_113_283 ();
 FILLCELL_X4 FILLER_0_113_295 ();
 FILLCELL_X1 FILLER_0_113_309 ();
 FILLCELL_X2 FILLER_0_113_324 ();
 FILLCELL_X4 FILLER_0_113_356 ();
 FILLCELL_X1 FILLER_0_113_360 ();
 FILLCELL_X1 FILLER_0_113_406 ();
 FILLCELL_X8 FILLER_0_113_421 ();
 FILLCELL_X2 FILLER_0_113_429 ();
 FILLCELL_X2 FILLER_0_113_438 ();
 FILLCELL_X1 FILLER_0_113_440 ();
 FILLCELL_X4 FILLER_0_113_466 ();
 FILLCELL_X1 FILLER_0_113_490 ();
 FILLCELL_X1 FILLER_0_113_506 ();
 FILLCELL_X1 FILLER_0_113_522 ();
 FILLCELL_X2 FILLER_0_113_537 ();
 FILLCELL_X1 FILLER_0_113_539 ();
 FILLCELL_X2 FILLER_0_113_550 ();
 FILLCELL_X2 FILLER_0_113_556 ();
 FILLCELL_X1 FILLER_0_113_558 ();
 FILLCELL_X2 FILLER_0_113_569 ();
 FILLCELL_X1 FILLER_0_113_571 ();
 FILLCELL_X8 FILLER_0_113_591 ();
 FILLCELL_X4 FILLER_0_113_599 ();
 FILLCELL_X2 FILLER_0_113_603 ();
 FILLCELL_X1 FILLER_0_113_605 ();
 FILLCELL_X8 FILLER_0_113_641 ();
 FILLCELL_X1 FILLER_0_113_659 ();
 FILLCELL_X1 FILLER_0_113_669 ();
 FILLCELL_X1 FILLER_0_113_680 ();
 FILLCELL_X1 FILLER_0_113_686 ();
 FILLCELL_X2 FILLER_0_113_696 ();
 FILLCELL_X4 FILLER_0_113_718 ();
 FILLCELL_X2 FILLER_0_113_727 ();
 FILLCELL_X1 FILLER_0_113_729 ();
 FILLCELL_X2 FILLER_0_113_740 ();
 FILLCELL_X4 FILLER_0_113_762 ();
 FILLCELL_X2 FILLER_0_113_766 ();
 FILLCELL_X8 FILLER_0_113_778 ();
 FILLCELL_X2 FILLER_0_113_786 ();
 FILLCELL_X16 FILLER_0_113_803 ();
 FILLCELL_X4 FILLER_0_113_819 ();
 FILLCELL_X1 FILLER_0_113_823 ();
 FILLCELL_X4 FILLER_0_113_849 ();
 FILLCELL_X8 FILLER_0_113_863 ();
 FILLCELL_X2 FILLER_0_113_871 ();
 FILLCELL_X8 FILLER_0_113_880 ();
 FILLCELL_X2 FILLER_0_113_888 ();
 FILLCELL_X1 FILLER_0_113_900 ();
 FILLCELL_X1 FILLER_0_113_925 ();
 FILLCELL_X4 FILLER_0_113_933 ();
 FILLCELL_X4 FILLER_0_113_969 ();
 FILLCELL_X2 FILLER_0_113_993 ();
 FILLCELL_X1 FILLER_0_113_995 ();
 FILLCELL_X32 FILLER_0_113_1010 ();
 FILLCELL_X32 FILLER_0_113_1042 ();
 FILLCELL_X32 FILLER_0_113_1074 ();
 FILLCELL_X32 FILLER_0_113_1106 ();
 FILLCELL_X8 FILLER_0_113_1138 ();
 FILLCELL_X2 FILLER_0_113_1146 ();
 FILLCELL_X32 FILLER_0_114_1 ();
 FILLCELL_X32 FILLER_0_114_33 ();
 FILLCELL_X32 FILLER_0_114_65 ();
 FILLCELL_X32 FILLER_0_114_97 ();
 FILLCELL_X32 FILLER_0_114_129 ();
 FILLCELL_X32 FILLER_0_114_161 ();
 FILLCELL_X32 FILLER_0_114_193 ();
 FILLCELL_X4 FILLER_0_114_225 ();
 FILLCELL_X1 FILLER_0_114_229 ();
 FILLCELL_X2 FILLER_0_114_250 ();
 FILLCELL_X2 FILLER_0_114_257 ();
 FILLCELL_X2 FILLER_0_114_279 ();
 FILLCELL_X1 FILLER_0_114_281 ();
 FILLCELL_X4 FILLER_0_114_297 ();
 FILLCELL_X2 FILLER_0_114_355 ();
 FILLCELL_X16 FILLER_0_114_367 ();
 FILLCELL_X4 FILLER_0_114_383 ();
 FILLCELL_X2 FILLER_0_114_387 ();
 FILLCELL_X32 FILLER_0_114_404 ();
 FILLCELL_X8 FILLER_0_114_436 ();
 FILLCELL_X2 FILLER_0_114_454 ();
 FILLCELL_X8 FILLER_0_114_465 ();
 FILLCELL_X2 FILLER_0_114_473 ();
 FILLCELL_X1 FILLER_0_114_475 ();
 FILLCELL_X1 FILLER_0_114_491 ();
 FILLCELL_X1 FILLER_0_114_502 ();
 FILLCELL_X2 FILLER_0_114_523 ();
 FILLCELL_X1 FILLER_0_114_525 ();
 FILLCELL_X2 FILLER_0_114_531 ();
 FILLCELL_X1 FILLER_0_114_562 ();
 FILLCELL_X1 FILLER_0_114_588 ();
 FILLCELL_X2 FILLER_0_114_599 ();
 FILLCELL_X2 FILLER_0_114_619 ();
 FILLCELL_X16 FILLER_0_114_632 ();
 FILLCELL_X4 FILLER_0_114_648 ();
 FILLCELL_X1 FILLER_0_114_667 ();
 FILLCELL_X1 FILLER_0_114_677 ();
 FILLCELL_X2 FILLER_0_114_688 ();
 FILLCELL_X1 FILLER_0_114_695 ();
 FILLCELL_X2 FILLER_0_114_706 ();
 FILLCELL_X1 FILLER_0_114_751 ();
 FILLCELL_X2 FILLER_0_114_781 ();
 FILLCELL_X1 FILLER_0_114_783 ();
 FILLCELL_X4 FILLER_0_114_802 ();
 FILLCELL_X1 FILLER_0_114_806 ();
 FILLCELL_X8 FILLER_0_114_817 ();
 FILLCELL_X4 FILLER_0_114_825 ();
 FILLCELL_X2 FILLER_0_114_829 ();
 FILLCELL_X32 FILLER_0_114_856 ();
 FILLCELL_X4 FILLER_0_114_888 ();
 FILLCELL_X8 FILLER_0_114_902 ();
 FILLCELL_X1 FILLER_0_114_910 ();
 FILLCELL_X2 FILLER_0_114_931 ();
 FILLCELL_X1 FILLER_0_114_933 ();
 FILLCELL_X2 FILLER_0_114_944 ();
 FILLCELL_X1 FILLER_0_114_946 ();
 FILLCELL_X2 FILLER_0_114_964 ();
 FILLCELL_X2 FILLER_0_114_976 ();
 FILLCELL_X32 FILLER_0_114_1008 ();
 FILLCELL_X32 FILLER_0_114_1040 ();
 FILLCELL_X32 FILLER_0_114_1072 ();
 FILLCELL_X32 FILLER_0_114_1104 ();
 FILLCELL_X8 FILLER_0_114_1136 ();
 FILLCELL_X4 FILLER_0_114_1144 ();
 FILLCELL_X32 FILLER_0_115_1 ();
 FILLCELL_X32 FILLER_0_115_33 ();
 FILLCELL_X32 FILLER_0_115_65 ();
 FILLCELL_X32 FILLER_0_115_97 ();
 FILLCELL_X32 FILLER_0_115_129 ();
 FILLCELL_X32 FILLER_0_115_161 ();
 FILLCELL_X32 FILLER_0_115_193 ();
 FILLCELL_X32 FILLER_0_115_225 ();
 FILLCELL_X16 FILLER_0_115_257 ();
 FILLCELL_X2 FILLER_0_115_273 ();
 FILLCELL_X1 FILLER_0_115_275 ();
 FILLCELL_X32 FILLER_0_115_286 ();
 FILLCELL_X2 FILLER_0_115_318 ();
 FILLCELL_X32 FILLER_0_115_335 ();
 FILLCELL_X32 FILLER_0_115_367 ();
 FILLCELL_X32 FILLER_0_115_399 ();
 FILLCELL_X8 FILLER_0_115_431 ();
 FILLCELL_X2 FILLER_0_115_439 ();
 FILLCELL_X1 FILLER_0_115_441 ();
 FILLCELL_X1 FILLER_0_115_467 ();
 FILLCELL_X4 FILLER_0_115_478 ();
 FILLCELL_X2 FILLER_0_115_482 ();
 FILLCELL_X2 FILLER_0_115_499 ();
 FILLCELL_X1 FILLER_0_115_501 ();
 FILLCELL_X1 FILLER_0_115_507 ();
 FILLCELL_X2 FILLER_0_115_563 ();
 FILLCELL_X8 FILLER_0_115_574 ();
 FILLCELL_X2 FILLER_0_115_582 ();
 FILLCELL_X1 FILLER_0_115_584 ();
 FILLCELL_X1 FILLER_0_115_590 ();
 FILLCELL_X2 FILLER_0_115_601 ();
 FILLCELL_X1 FILLER_0_115_603 ();
 FILLCELL_X16 FILLER_0_115_624 ();
 FILLCELL_X8 FILLER_0_115_640 ();
 FILLCELL_X4 FILLER_0_115_648 ();
 FILLCELL_X4 FILLER_0_115_662 ();
 FILLCELL_X2 FILLER_0_115_666 ();
 FILLCELL_X1 FILLER_0_115_668 ();
 FILLCELL_X2 FILLER_0_115_699 ();
 FILLCELL_X1 FILLER_0_115_721 ();
 FILLCELL_X2 FILLER_0_115_732 ();
 FILLCELL_X1 FILLER_0_115_744 ();
 FILLCELL_X2 FILLER_0_115_765 ();
 FILLCELL_X1 FILLER_0_115_767 ();
 FILLCELL_X4 FILLER_0_115_773 ();
 FILLCELL_X4 FILLER_0_115_782 ();
 FILLCELL_X32 FILLER_0_115_820 ();
 FILLCELL_X4 FILLER_0_115_852 ();
 FILLCELL_X4 FILLER_0_115_866 ();
 FILLCELL_X2 FILLER_0_115_870 ();
 FILLCELL_X4 FILLER_0_115_882 ();
 FILLCELL_X1 FILLER_0_115_886 ();
 FILLCELL_X1 FILLER_0_115_922 ();
 FILLCELL_X4 FILLER_0_115_943 ();
 FILLCELL_X2 FILLER_0_115_947 ();
 FILLCELL_X1 FILLER_0_115_959 ();
 FILLCELL_X2 FILLER_0_115_985 ();
 FILLCELL_X32 FILLER_0_115_1001 ();
 FILLCELL_X32 FILLER_0_115_1033 ();
 FILLCELL_X32 FILLER_0_115_1065 ();
 FILLCELL_X32 FILLER_0_115_1097 ();
 FILLCELL_X16 FILLER_0_115_1129 ();
 FILLCELL_X2 FILLER_0_115_1145 ();
 FILLCELL_X1 FILLER_0_115_1147 ();
 FILLCELL_X32 FILLER_0_116_1 ();
 FILLCELL_X32 FILLER_0_116_33 ();
 FILLCELL_X32 FILLER_0_116_65 ();
 FILLCELL_X32 FILLER_0_116_97 ();
 FILLCELL_X32 FILLER_0_116_129 ();
 FILLCELL_X32 FILLER_0_116_161 ();
 FILLCELL_X32 FILLER_0_116_193 ();
 FILLCELL_X32 FILLER_0_116_225 ();
 FILLCELL_X32 FILLER_0_116_257 ();
 FILLCELL_X32 FILLER_0_116_289 ();
 FILLCELL_X32 FILLER_0_116_321 ();
 FILLCELL_X32 FILLER_0_116_353 ();
 FILLCELL_X32 FILLER_0_116_385 ();
 FILLCELL_X32 FILLER_0_116_417 ();
 FILLCELL_X16 FILLER_0_116_449 ();
 FILLCELL_X1 FILLER_0_116_465 ();
 FILLCELL_X2 FILLER_0_116_505 ();
 FILLCELL_X1 FILLER_0_116_507 ();
 FILLCELL_X2 FILLER_0_116_538 ();
 FILLCELL_X2 FILLER_0_116_560 ();
 FILLCELL_X4 FILLER_0_116_592 ();
 FILLCELL_X1 FILLER_0_116_596 ();
 FILLCELL_X16 FILLER_0_116_607 ();
 FILLCELL_X8 FILLER_0_116_623 ();
 FILLCELL_X16 FILLER_0_116_632 ();
 FILLCELL_X8 FILLER_0_116_648 ();
 FILLCELL_X4 FILLER_0_116_656 ();
 FILLCELL_X2 FILLER_0_116_660 ();
 FILLCELL_X1 FILLER_0_116_681 ();
 FILLCELL_X1 FILLER_0_116_692 ();
 FILLCELL_X1 FILLER_0_116_703 ();
 FILLCELL_X1 FILLER_0_116_714 ();
 FILLCELL_X2 FILLER_0_116_720 ();
 FILLCELL_X1 FILLER_0_116_722 ();
 FILLCELL_X1 FILLER_0_116_733 ();
 FILLCELL_X1 FILLER_0_116_784 ();
 FILLCELL_X16 FILLER_0_116_815 ();
 FILLCELL_X8 FILLER_0_116_831 ();
 FILLCELL_X4 FILLER_0_116_839 ();
 FILLCELL_X2 FILLER_0_116_983 ();
 FILLCELL_X32 FILLER_0_116_1005 ();
 FILLCELL_X32 FILLER_0_116_1037 ();
 FILLCELL_X32 FILLER_0_116_1069 ();
 FILLCELL_X32 FILLER_0_116_1101 ();
 FILLCELL_X8 FILLER_0_116_1133 ();
 FILLCELL_X4 FILLER_0_116_1141 ();
 FILLCELL_X2 FILLER_0_116_1145 ();
 FILLCELL_X1 FILLER_0_116_1147 ();
 FILLCELL_X32 FILLER_0_117_1 ();
 FILLCELL_X32 FILLER_0_117_33 ();
 FILLCELL_X32 FILLER_0_117_65 ();
 FILLCELL_X32 FILLER_0_117_97 ();
 FILLCELL_X32 FILLER_0_117_129 ();
 FILLCELL_X32 FILLER_0_117_161 ();
 FILLCELL_X32 FILLER_0_117_193 ();
 FILLCELL_X32 FILLER_0_117_225 ();
 FILLCELL_X32 FILLER_0_117_257 ();
 FILLCELL_X32 FILLER_0_117_289 ();
 FILLCELL_X32 FILLER_0_117_321 ();
 FILLCELL_X32 FILLER_0_117_353 ();
 FILLCELL_X32 FILLER_0_117_385 ();
 FILLCELL_X32 FILLER_0_117_417 ();
 FILLCELL_X2 FILLER_0_117_449 ();
 FILLCELL_X1 FILLER_0_117_451 ();
 FILLCELL_X32 FILLER_0_117_462 ();
 FILLCELL_X8 FILLER_0_117_494 ();
 FILLCELL_X16 FILLER_0_117_512 ();
 FILLCELL_X8 FILLER_0_117_528 ();
 FILLCELL_X2 FILLER_0_117_536 ();
 FILLCELL_X1 FILLER_0_117_538 ();
 FILLCELL_X8 FILLER_0_117_549 ();
 FILLCELL_X4 FILLER_0_117_557 ();
 FILLCELL_X1 FILLER_0_117_561 ();
 FILLCELL_X32 FILLER_0_117_572 ();
 FILLCELL_X32 FILLER_0_117_604 ();
 FILLCELL_X32 FILLER_0_117_636 ();
 FILLCELL_X16 FILLER_0_117_668 ();
 FILLCELL_X1 FILLER_0_117_684 ();
 FILLCELL_X16 FILLER_0_117_695 ();
 FILLCELL_X4 FILLER_0_117_711 ();
 FILLCELL_X2 FILLER_0_117_715 ();
 FILLCELL_X1 FILLER_0_117_727 ();
 FILLCELL_X1 FILLER_0_117_738 ();
 FILLCELL_X1 FILLER_0_117_744 ();
 FILLCELL_X1 FILLER_0_117_755 ();
 FILLCELL_X4 FILLER_0_117_761 ();
 FILLCELL_X32 FILLER_0_117_775 ();
 FILLCELL_X32 FILLER_0_117_807 ();
 FILLCELL_X8 FILLER_0_117_839 ();
 FILLCELL_X4 FILLER_0_117_847 ();
 FILLCELL_X1 FILLER_0_117_851 ();
 FILLCELL_X4 FILLER_0_117_872 ();
 FILLCELL_X1 FILLER_0_117_876 ();
 FILLCELL_X1 FILLER_0_117_882 ();
 FILLCELL_X1 FILLER_0_117_898 ();
 FILLCELL_X1 FILLER_0_117_904 ();
 FILLCELL_X2 FILLER_0_117_910 ();
 FILLCELL_X1 FILLER_0_117_912 ();
 FILLCELL_X2 FILLER_0_117_923 ();
 FILLCELL_X2 FILLER_0_117_935 ();
 FILLCELL_X1 FILLER_0_117_937 ();
 FILLCELL_X4 FILLER_0_117_963 ();
 FILLCELL_X32 FILLER_0_117_977 ();
 FILLCELL_X32 FILLER_0_117_1009 ();
 FILLCELL_X32 FILLER_0_117_1041 ();
 FILLCELL_X32 FILLER_0_117_1073 ();
 FILLCELL_X32 FILLER_0_117_1105 ();
 FILLCELL_X8 FILLER_0_117_1137 ();
 FILLCELL_X2 FILLER_0_117_1145 ();
 FILLCELL_X1 FILLER_0_117_1147 ();
 FILLCELL_X32 FILLER_0_118_1 ();
 FILLCELL_X32 FILLER_0_118_33 ();
 FILLCELL_X32 FILLER_0_118_65 ();
 FILLCELL_X32 FILLER_0_118_97 ();
 FILLCELL_X32 FILLER_0_118_129 ();
 FILLCELL_X32 FILLER_0_118_161 ();
 FILLCELL_X32 FILLER_0_118_193 ();
 FILLCELL_X32 FILLER_0_118_225 ();
 FILLCELL_X32 FILLER_0_118_257 ();
 FILLCELL_X32 FILLER_0_118_289 ();
 FILLCELL_X32 FILLER_0_118_321 ();
 FILLCELL_X32 FILLER_0_118_353 ();
 FILLCELL_X32 FILLER_0_118_385 ();
 FILLCELL_X32 FILLER_0_118_417 ();
 FILLCELL_X32 FILLER_0_118_449 ();
 FILLCELL_X32 FILLER_0_118_481 ();
 FILLCELL_X32 FILLER_0_118_513 ();
 FILLCELL_X32 FILLER_0_118_545 ();
 FILLCELL_X32 FILLER_0_118_577 ();
 FILLCELL_X16 FILLER_0_118_609 ();
 FILLCELL_X4 FILLER_0_118_625 ();
 FILLCELL_X2 FILLER_0_118_629 ();
 FILLCELL_X32 FILLER_0_118_632 ();
 FILLCELL_X32 FILLER_0_118_664 ();
 FILLCELL_X32 FILLER_0_118_696 ();
 FILLCELL_X16 FILLER_0_118_728 ();
 FILLCELL_X4 FILLER_0_118_744 ();
 FILLCELL_X2 FILLER_0_118_748 ();
 FILLCELL_X32 FILLER_0_118_760 ();
 FILLCELL_X32 FILLER_0_118_792 ();
 FILLCELL_X32 FILLER_0_118_824 ();
 FILLCELL_X16 FILLER_0_118_856 ();
 FILLCELL_X8 FILLER_0_118_872 ();
 FILLCELL_X2 FILLER_0_118_880 ();
 FILLCELL_X1 FILLER_0_118_882 ();
 FILLCELL_X8 FILLER_0_118_893 ();
 FILLCELL_X2 FILLER_0_118_901 ();
 FILLCELL_X8 FILLER_0_118_913 ();
 FILLCELL_X4 FILLER_0_118_921 ();
 FILLCELL_X1 FILLER_0_118_925 ();
 FILLCELL_X16 FILLER_0_118_936 ();
 FILLCELL_X8 FILLER_0_118_952 ();
 FILLCELL_X2 FILLER_0_118_960 ();
 FILLCELL_X32 FILLER_0_118_967 ();
 FILLCELL_X32 FILLER_0_118_999 ();
 FILLCELL_X32 FILLER_0_118_1031 ();
 FILLCELL_X32 FILLER_0_118_1063 ();
 FILLCELL_X32 FILLER_0_118_1095 ();
 FILLCELL_X16 FILLER_0_118_1127 ();
 FILLCELL_X4 FILLER_0_118_1143 ();
 FILLCELL_X1 FILLER_0_118_1147 ();
 FILLCELL_X32 FILLER_0_119_1 ();
 FILLCELL_X32 FILLER_0_119_33 ();
 FILLCELL_X32 FILLER_0_119_65 ();
 FILLCELL_X32 FILLER_0_119_97 ();
 FILLCELL_X32 FILLER_0_119_129 ();
 FILLCELL_X32 FILLER_0_119_161 ();
 FILLCELL_X32 FILLER_0_119_193 ();
 FILLCELL_X32 FILLER_0_119_225 ();
 FILLCELL_X32 FILLER_0_119_257 ();
 FILLCELL_X32 FILLER_0_119_289 ();
 FILLCELL_X32 FILLER_0_119_321 ();
 FILLCELL_X32 FILLER_0_119_353 ();
 FILLCELL_X32 FILLER_0_119_385 ();
 FILLCELL_X32 FILLER_0_119_417 ();
 FILLCELL_X32 FILLER_0_119_449 ();
 FILLCELL_X32 FILLER_0_119_481 ();
 FILLCELL_X32 FILLER_0_119_513 ();
 FILLCELL_X32 FILLER_0_119_545 ();
 FILLCELL_X32 FILLER_0_119_577 ();
 FILLCELL_X32 FILLER_0_119_609 ();
 FILLCELL_X32 FILLER_0_119_641 ();
 FILLCELL_X32 FILLER_0_119_673 ();
 FILLCELL_X32 FILLER_0_119_705 ();
 FILLCELL_X32 FILLER_0_119_737 ();
 FILLCELL_X32 FILLER_0_119_769 ();
 FILLCELL_X32 FILLER_0_119_801 ();
 FILLCELL_X32 FILLER_0_119_833 ();
 FILLCELL_X32 FILLER_0_119_865 ();
 FILLCELL_X32 FILLER_0_119_897 ();
 FILLCELL_X32 FILLER_0_119_929 ();
 FILLCELL_X32 FILLER_0_119_961 ();
 FILLCELL_X32 FILLER_0_119_993 ();
 FILLCELL_X32 FILLER_0_119_1025 ();
 FILLCELL_X32 FILLER_0_119_1057 ();
 FILLCELL_X32 FILLER_0_119_1089 ();
 FILLCELL_X16 FILLER_0_119_1121 ();
 FILLCELL_X8 FILLER_0_119_1137 ();
 FILLCELL_X2 FILLER_0_119_1145 ();
 FILLCELL_X1 FILLER_0_119_1147 ();
 FILLCELL_X32 FILLER_0_120_1 ();
 FILLCELL_X32 FILLER_0_120_33 ();
 FILLCELL_X32 FILLER_0_120_65 ();
 FILLCELL_X32 FILLER_0_120_97 ();
 FILLCELL_X32 FILLER_0_120_129 ();
 FILLCELL_X32 FILLER_0_120_161 ();
 FILLCELL_X32 FILLER_0_120_193 ();
 FILLCELL_X32 FILLER_0_120_225 ();
 FILLCELL_X32 FILLER_0_120_257 ();
 FILLCELL_X32 FILLER_0_120_289 ();
 FILLCELL_X32 FILLER_0_120_321 ();
 FILLCELL_X32 FILLER_0_120_353 ();
 FILLCELL_X32 FILLER_0_120_385 ();
 FILLCELL_X32 FILLER_0_120_417 ();
 FILLCELL_X32 FILLER_0_120_449 ();
 FILLCELL_X32 FILLER_0_120_481 ();
 FILLCELL_X32 FILLER_0_120_513 ();
 FILLCELL_X32 FILLER_0_120_545 ();
 FILLCELL_X32 FILLER_0_120_577 ();
 FILLCELL_X16 FILLER_0_120_609 ();
 FILLCELL_X4 FILLER_0_120_625 ();
 FILLCELL_X2 FILLER_0_120_629 ();
 FILLCELL_X32 FILLER_0_120_632 ();
 FILLCELL_X32 FILLER_0_120_664 ();
 FILLCELL_X32 FILLER_0_120_696 ();
 FILLCELL_X32 FILLER_0_120_728 ();
 FILLCELL_X32 FILLER_0_120_760 ();
 FILLCELL_X32 FILLER_0_120_792 ();
 FILLCELL_X32 FILLER_0_120_824 ();
 FILLCELL_X32 FILLER_0_120_856 ();
 FILLCELL_X32 FILLER_0_120_888 ();
 FILLCELL_X32 FILLER_0_120_920 ();
 FILLCELL_X32 FILLER_0_120_952 ();
 FILLCELL_X32 FILLER_0_120_984 ();
 FILLCELL_X32 FILLER_0_120_1016 ();
 FILLCELL_X32 FILLER_0_120_1048 ();
 FILLCELL_X32 FILLER_0_120_1080 ();
 FILLCELL_X32 FILLER_0_120_1112 ();
 FILLCELL_X4 FILLER_0_120_1144 ();
 FILLCELL_X32 FILLER_0_121_1 ();
 FILLCELL_X32 FILLER_0_121_33 ();
 FILLCELL_X32 FILLER_0_121_65 ();
 FILLCELL_X32 FILLER_0_121_97 ();
 FILLCELL_X32 FILLER_0_121_129 ();
 FILLCELL_X32 FILLER_0_121_161 ();
 FILLCELL_X32 FILLER_0_121_193 ();
 FILLCELL_X32 FILLER_0_121_225 ();
 FILLCELL_X32 FILLER_0_121_257 ();
 FILLCELL_X32 FILLER_0_121_289 ();
 FILLCELL_X32 FILLER_0_121_321 ();
 FILLCELL_X32 FILLER_0_121_353 ();
 FILLCELL_X32 FILLER_0_121_385 ();
 FILLCELL_X32 FILLER_0_121_417 ();
 FILLCELL_X32 FILLER_0_121_449 ();
 FILLCELL_X32 FILLER_0_121_481 ();
 FILLCELL_X32 FILLER_0_121_513 ();
 FILLCELL_X32 FILLER_0_121_545 ();
 FILLCELL_X32 FILLER_0_121_577 ();
 FILLCELL_X32 FILLER_0_121_609 ();
 FILLCELL_X32 FILLER_0_121_641 ();
 FILLCELL_X32 FILLER_0_121_673 ();
 FILLCELL_X32 FILLER_0_121_705 ();
 FILLCELL_X32 FILLER_0_121_737 ();
 FILLCELL_X32 FILLER_0_121_769 ();
 FILLCELL_X32 FILLER_0_121_801 ();
 FILLCELL_X32 FILLER_0_121_833 ();
 FILLCELL_X32 FILLER_0_121_865 ();
 FILLCELL_X32 FILLER_0_121_897 ();
 FILLCELL_X32 FILLER_0_121_929 ();
 FILLCELL_X32 FILLER_0_121_961 ();
 FILLCELL_X32 FILLER_0_121_993 ();
 FILLCELL_X32 FILLER_0_121_1025 ();
 FILLCELL_X32 FILLER_0_121_1057 ();
 FILLCELL_X32 FILLER_0_121_1089 ();
 FILLCELL_X16 FILLER_0_121_1121 ();
 FILLCELL_X8 FILLER_0_121_1137 ();
 FILLCELL_X2 FILLER_0_121_1145 ();
 FILLCELL_X1 FILLER_0_121_1147 ();
 FILLCELL_X32 FILLER_0_122_1 ();
 FILLCELL_X32 FILLER_0_122_33 ();
 FILLCELL_X32 FILLER_0_122_65 ();
 FILLCELL_X32 FILLER_0_122_97 ();
 FILLCELL_X32 FILLER_0_122_129 ();
 FILLCELL_X32 FILLER_0_122_161 ();
 FILLCELL_X32 FILLER_0_122_193 ();
 FILLCELL_X32 FILLER_0_122_225 ();
 FILLCELL_X32 FILLER_0_122_257 ();
 FILLCELL_X32 FILLER_0_122_289 ();
 FILLCELL_X32 FILLER_0_122_321 ();
 FILLCELL_X32 FILLER_0_122_353 ();
 FILLCELL_X32 FILLER_0_122_385 ();
 FILLCELL_X32 FILLER_0_122_417 ();
 FILLCELL_X32 FILLER_0_122_449 ();
 FILLCELL_X32 FILLER_0_122_481 ();
 FILLCELL_X32 FILLER_0_122_513 ();
 FILLCELL_X32 FILLER_0_122_545 ();
 FILLCELL_X32 FILLER_0_122_577 ();
 FILLCELL_X16 FILLER_0_122_609 ();
 FILLCELL_X4 FILLER_0_122_625 ();
 FILLCELL_X2 FILLER_0_122_629 ();
 FILLCELL_X32 FILLER_0_122_632 ();
 FILLCELL_X32 FILLER_0_122_664 ();
 FILLCELL_X32 FILLER_0_122_696 ();
 FILLCELL_X32 FILLER_0_122_728 ();
 FILLCELL_X32 FILLER_0_122_760 ();
 FILLCELL_X32 FILLER_0_122_792 ();
 FILLCELL_X32 FILLER_0_122_824 ();
 FILLCELL_X32 FILLER_0_122_856 ();
 FILLCELL_X32 FILLER_0_122_888 ();
 FILLCELL_X32 FILLER_0_122_920 ();
 FILLCELL_X32 FILLER_0_122_952 ();
 FILLCELL_X32 FILLER_0_122_984 ();
 FILLCELL_X32 FILLER_0_122_1016 ();
 FILLCELL_X32 FILLER_0_122_1048 ();
 FILLCELL_X32 FILLER_0_122_1080 ();
 FILLCELL_X32 FILLER_0_122_1112 ();
 FILLCELL_X4 FILLER_0_122_1144 ();
 FILLCELL_X32 FILLER_0_123_1 ();
 FILLCELL_X32 FILLER_0_123_33 ();
 FILLCELL_X32 FILLER_0_123_65 ();
 FILLCELL_X32 FILLER_0_123_97 ();
 FILLCELL_X32 FILLER_0_123_129 ();
 FILLCELL_X32 FILLER_0_123_161 ();
 FILLCELL_X32 FILLER_0_123_193 ();
 FILLCELL_X32 FILLER_0_123_225 ();
 FILLCELL_X32 FILLER_0_123_257 ();
 FILLCELL_X32 FILLER_0_123_289 ();
 FILLCELL_X32 FILLER_0_123_321 ();
 FILLCELL_X32 FILLER_0_123_353 ();
 FILLCELL_X32 FILLER_0_123_385 ();
 FILLCELL_X32 FILLER_0_123_417 ();
 FILLCELL_X32 FILLER_0_123_449 ();
 FILLCELL_X32 FILLER_0_123_481 ();
 FILLCELL_X32 FILLER_0_123_513 ();
 FILLCELL_X32 FILLER_0_123_545 ();
 FILLCELL_X32 FILLER_0_123_577 ();
 FILLCELL_X32 FILLER_0_123_609 ();
 FILLCELL_X32 FILLER_0_123_641 ();
 FILLCELL_X32 FILLER_0_123_673 ();
 FILLCELL_X32 FILLER_0_123_705 ();
 FILLCELL_X32 FILLER_0_123_737 ();
 FILLCELL_X32 FILLER_0_123_769 ();
 FILLCELL_X32 FILLER_0_123_801 ();
 FILLCELL_X32 FILLER_0_123_833 ();
 FILLCELL_X32 FILLER_0_123_865 ();
 FILLCELL_X32 FILLER_0_123_897 ();
 FILLCELL_X32 FILLER_0_123_929 ();
 FILLCELL_X32 FILLER_0_123_961 ();
 FILLCELL_X32 FILLER_0_123_993 ();
 FILLCELL_X32 FILLER_0_123_1025 ();
 FILLCELL_X32 FILLER_0_123_1057 ();
 FILLCELL_X32 FILLER_0_123_1089 ();
 FILLCELL_X16 FILLER_0_123_1121 ();
 FILLCELL_X8 FILLER_0_123_1137 ();
 FILLCELL_X2 FILLER_0_123_1145 ();
 FILLCELL_X1 FILLER_0_123_1147 ();
 FILLCELL_X32 FILLER_0_124_1 ();
 FILLCELL_X32 FILLER_0_124_33 ();
 FILLCELL_X32 FILLER_0_124_65 ();
 FILLCELL_X32 FILLER_0_124_97 ();
 FILLCELL_X32 FILLER_0_124_129 ();
 FILLCELL_X32 FILLER_0_124_161 ();
 FILLCELL_X32 FILLER_0_124_193 ();
 FILLCELL_X32 FILLER_0_124_225 ();
 FILLCELL_X32 FILLER_0_124_257 ();
 FILLCELL_X32 FILLER_0_124_289 ();
 FILLCELL_X32 FILLER_0_124_321 ();
 FILLCELL_X32 FILLER_0_124_353 ();
 FILLCELL_X32 FILLER_0_124_385 ();
 FILLCELL_X32 FILLER_0_124_417 ();
 FILLCELL_X32 FILLER_0_124_449 ();
 FILLCELL_X32 FILLER_0_124_481 ();
 FILLCELL_X32 FILLER_0_124_513 ();
 FILLCELL_X32 FILLER_0_124_545 ();
 FILLCELL_X32 FILLER_0_124_577 ();
 FILLCELL_X16 FILLER_0_124_609 ();
 FILLCELL_X4 FILLER_0_124_625 ();
 FILLCELL_X2 FILLER_0_124_629 ();
 FILLCELL_X32 FILLER_0_124_632 ();
 FILLCELL_X32 FILLER_0_124_664 ();
 FILLCELL_X32 FILLER_0_124_696 ();
 FILLCELL_X32 FILLER_0_124_728 ();
 FILLCELL_X32 FILLER_0_124_760 ();
 FILLCELL_X32 FILLER_0_124_792 ();
 FILLCELL_X32 FILLER_0_124_824 ();
 FILLCELL_X32 FILLER_0_124_856 ();
 FILLCELL_X32 FILLER_0_124_888 ();
 FILLCELL_X32 FILLER_0_124_920 ();
 FILLCELL_X32 FILLER_0_124_952 ();
 FILLCELL_X32 FILLER_0_124_984 ();
 FILLCELL_X32 FILLER_0_124_1016 ();
 FILLCELL_X32 FILLER_0_124_1048 ();
 FILLCELL_X32 FILLER_0_124_1080 ();
 FILLCELL_X32 FILLER_0_124_1112 ();
 FILLCELL_X4 FILLER_0_124_1144 ();
 FILLCELL_X32 FILLER_0_125_1 ();
 FILLCELL_X32 FILLER_0_125_33 ();
 FILLCELL_X32 FILLER_0_125_65 ();
 FILLCELL_X32 FILLER_0_125_97 ();
 FILLCELL_X32 FILLER_0_125_129 ();
 FILLCELL_X32 FILLER_0_125_161 ();
 FILLCELL_X32 FILLER_0_125_193 ();
 FILLCELL_X32 FILLER_0_125_225 ();
 FILLCELL_X32 FILLER_0_125_257 ();
 FILLCELL_X32 FILLER_0_125_289 ();
 FILLCELL_X32 FILLER_0_125_321 ();
 FILLCELL_X32 FILLER_0_125_353 ();
 FILLCELL_X32 FILLER_0_125_385 ();
 FILLCELL_X32 FILLER_0_125_417 ();
 FILLCELL_X32 FILLER_0_125_449 ();
 FILLCELL_X32 FILLER_0_125_481 ();
 FILLCELL_X32 FILLER_0_125_513 ();
 FILLCELL_X32 FILLER_0_125_545 ();
 FILLCELL_X32 FILLER_0_125_577 ();
 FILLCELL_X32 FILLER_0_125_609 ();
 FILLCELL_X32 FILLER_0_125_641 ();
 FILLCELL_X32 FILLER_0_125_673 ();
 FILLCELL_X32 FILLER_0_125_705 ();
 FILLCELL_X32 FILLER_0_125_737 ();
 FILLCELL_X32 FILLER_0_125_769 ();
 FILLCELL_X32 FILLER_0_125_801 ();
 FILLCELL_X32 FILLER_0_125_833 ();
 FILLCELL_X32 FILLER_0_125_865 ();
 FILLCELL_X32 FILLER_0_125_897 ();
 FILLCELL_X32 FILLER_0_125_929 ();
 FILLCELL_X32 FILLER_0_125_961 ();
 FILLCELL_X32 FILLER_0_125_993 ();
 FILLCELL_X32 FILLER_0_125_1025 ();
 FILLCELL_X32 FILLER_0_125_1057 ();
 FILLCELL_X32 FILLER_0_125_1089 ();
 FILLCELL_X16 FILLER_0_125_1121 ();
 FILLCELL_X8 FILLER_0_125_1137 ();
 FILLCELL_X2 FILLER_0_125_1145 ();
 FILLCELL_X1 FILLER_0_125_1147 ();
 FILLCELL_X32 FILLER_0_126_1 ();
 FILLCELL_X32 FILLER_0_126_33 ();
 FILLCELL_X32 FILLER_0_126_65 ();
 FILLCELL_X32 FILLER_0_126_97 ();
 FILLCELL_X32 FILLER_0_126_129 ();
 FILLCELL_X32 FILLER_0_126_161 ();
 FILLCELL_X32 FILLER_0_126_193 ();
 FILLCELL_X32 FILLER_0_126_225 ();
 FILLCELL_X32 FILLER_0_126_257 ();
 FILLCELL_X32 FILLER_0_126_289 ();
 FILLCELL_X32 FILLER_0_126_321 ();
 FILLCELL_X32 FILLER_0_126_353 ();
 FILLCELL_X32 FILLER_0_126_385 ();
 FILLCELL_X32 FILLER_0_126_417 ();
 FILLCELL_X32 FILLER_0_126_449 ();
 FILLCELL_X32 FILLER_0_126_481 ();
 FILLCELL_X32 FILLER_0_126_513 ();
 FILLCELL_X32 FILLER_0_126_545 ();
 FILLCELL_X32 FILLER_0_126_577 ();
 FILLCELL_X16 FILLER_0_126_609 ();
 FILLCELL_X4 FILLER_0_126_625 ();
 FILLCELL_X2 FILLER_0_126_629 ();
 FILLCELL_X32 FILLER_0_126_632 ();
 FILLCELL_X32 FILLER_0_126_664 ();
 FILLCELL_X32 FILLER_0_126_696 ();
 FILLCELL_X32 FILLER_0_126_728 ();
 FILLCELL_X32 FILLER_0_126_760 ();
 FILLCELL_X32 FILLER_0_126_792 ();
 FILLCELL_X32 FILLER_0_126_824 ();
 FILLCELL_X32 FILLER_0_126_856 ();
 FILLCELL_X32 FILLER_0_126_888 ();
 FILLCELL_X32 FILLER_0_126_920 ();
 FILLCELL_X32 FILLER_0_126_952 ();
 FILLCELL_X32 FILLER_0_126_984 ();
 FILLCELL_X32 FILLER_0_126_1016 ();
 FILLCELL_X32 FILLER_0_126_1048 ();
 FILLCELL_X32 FILLER_0_126_1080 ();
 FILLCELL_X32 FILLER_0_126_1112 ();
 FILLCELL_X4 FILLER_0_126_1144 ();
 FILLCELL_X32 FILLER_0_127_1 ();
 FILLCELL_X32 FILLER_0_127_33 ();
 FILLCELL_X32 FILLER_0_127_65 ();
 FILLCELL_X32 FILLER_0_127_97 ();
 FILLCELL_X32 FILLER_0_127_129 ();
 FILLCELL_X32 FILLER_0_127_161 ();
 FILLCELL_X32 FILLER_0_127_193 ();
 FILLCELL_X32 FILLER_0_127_225 ();
 FILLCELL_X32 FILLER_0_127_257 ();
 FILLCELL_X32 FILLER_0_127_289 ();
 FILLCELL_X32 FILLER_0_127_321 ();
 FILLCELL_X32 FILLER_0_127_353 ();
 FILLCELL_X32 FILLER_0_127_385 ();
 FILLCELL_X32 FILLER_0_127_417 ();
 FILLCELL_X32 FILLER_0_127_449 ();
 FILLCELL_X32 FILLER_0_127_481 ();
 FILLCELL_X32 FILLER_0_127_513 ();
 FILLCELL_X32 FILLER_0_127_545 ();
 FILLCELL_X32 FILLER_0_127_577 ();
 FILLCELL_X32 FILLER_0_127_609 ();
 FILLCELL_X32 FILLER_0_127_641 ();
 FILLCELL_X32 FILLER_0_127_673 ();
 FILLCELL_X32 FILLER_0_127_705 ();
 FILLCELL_X32 FILLER_0_127_737 ();
 FILLCELL_X32 FILLER_0_127_769 ();
 FILLCELL_X32 FILLER_0_127_801 ();
 FILLCELL_X32 FILLER_0_127_833 ();
 FILLCELL_X32 FILLER_0_127_865 ();
 FILLCELL_X32 FILLER_0_127_897 ();
 FILLCELL_X32 FILLER_0_127_929 ();
 FILLCELL_X32 FILLER_0_127_961 ();
 FILLCELL_X32 FILLER_0_127_993 ();
 FILLCELL_X32 FILLER_0_127_1025 ();
 FILLCELL_X32 FILLER_0_127_1057 ();
 FILLCELL_X32 FILLER_0_127_1089 ();
 FILLCELL_X16 FILLER_0_127_1121 ();
 FILLCELL_X8 FILLER_0_127_1137 ();
 FILLCELL_X2 FILLER_0_127_1145 ();
 FILLCELL_X1 FILLER_0_127_1147 ();
 FILLCELL_X32 FILLER_0_128_1 ();
 FILLCELL_X32 FILLER_0_128_33 ();
 FILLCELL_X32 FILLER_0_128_65 ();
 FILLCELL_X32 FILLER_0_128_97 ();
 FILLCELL_X32 FILLER_0_128_129 ();
 FILLCELL_X32 FILLER_0_128_161 ();
 FILLCELL_X32 FILLER_0_128_193 ();
 FILLCELL_X32 FILLER_0_128_225 ();
 FILLCELL_X32 FILLER_0_128_257 ();
 FILLCELL_X32 FILLER_0_128_289 ();
 FILLCELL_X32 FILLER_0_128_321 ();
 FILLCELL_X32 FILLER_0_128_353 ();
 FILLCELL_X32 FILLER_0_128_385 ();
 FILLCELL_X32 FILLER_0_128_417 ();
 FILLCELL_X32 FILLER_0_128_449 ();
 FILLCELL_X32 FILLER_0_128_481 ();
 FILLCELL_X32 FILLER_0_128_513 ();
 FILLCELL_X32 FILLER_0_128_545 ();
 FILLCELL_X32 FILLER_0_128_577 ();
 FILLCELL_X16 FILLER_0_128_609 ();
 FILLCELL_X4 FILLER_0_128_625 ();
 FILLCELL_X2 FILLER_0_128_629 ();
 FILLCELL_X32 FILLER_0_128_632 ();
 FILLCELL_X32 FILLER_0_128_664 ();
 FILLCELL_X32 FILLER_0_128_696 ();
 FILLCELL_X32 FILLER_0_128_728 ();
 FILLCELL_X32 FILLER_0_128_760 ();
 FILLCELL_X32 FILLER_0_128_792 ();
 FILLCELL_X32 FILLER_0_128_824 ();
 FILLCELL_X32 FILLER_0_128_856 ();
 FILLCELL_X32 FILLER_0_128_888 ();
 FILLCELL_X32 FILLER_0_128_920 ();
 FILLCELL_X32 FILLER_0_128_952 ();
 FILLCELL_X32 FILLER_0_128_984 ();
 FILLCELL_X32 FILLER_0_128_1016 ();
 FILLCELL_X32 FILLER_0_128_1048 ();
 FILLCELL_X32 FILLER_0_128_1080 ();
 FILLCELL_X32 FILLER_0_128_1112 ();
 FILLCELL_X4 FILLER_0_128_1144 ();
 FILLCELL_X32 FILLER_0_129_1 ();
 FILLCELL_X32 FILLER_0_129_33 ();
 FILLCELL_X32 FILLER_0_129_65 ();
 FILLCELL_X32 FILLER_0_129_97 ();
 FILLCELL_X32 FILLER_0_129_129 ();
 FILLCELL_X32 FILLER_0_129_161 ();
 FILLCELL_X32 FILLER_0_129_193 ();
 FILLCELL_X32 FILLER_0_129_225 ();
 FILLCELL_X32 FILLER_0_129_257 ();
 FILLCELL_X32 FILLER_0_129_289 ();
 FILLCELL_X32 FILLER_0_129_321 ();
 FILLCELL_X32 FILLER_0_129_353 ();
 FILLCELL_X32 FILLER_0_129_385 ();
 FILLCELL_X32 FILLER_0_129_417 ();
 FILLCELL_X32 FILLER_0_129_449 ();
 FILLCELL_X32 FILLER_0_129_481 ();
 FILLCELL_X32 FILLER_0_129_513 ();
 FILLCELL_X32 FILLER_0_129_545 ();
 FILLCELL_X32 FILLER_0_129_577 ();
 FILLCELL_X32 FILLER_0_129_609 ();
 FILLCELL_X32 FILLER_0_129_641 ();
 FILLCELL_X32 FILLER_0_129_673 ();
 FILLCELL_X32 FILLER_0_129_705 ();
 FILLCELL_X32 FILLER_0_129_737 ();
 FILLCELL_X32 FILLER_0_129_769 ();
 FILLCELL_X32 FILLER_0_129_801 ();
 FILLCELL_X32 FILLER_0_129_833 ();
 FILLCELL_X32 FILLER_0_129_865 ();
 FILLCELL_X32 FILLER_0_129_897 ();
 FILLCELL_X32 FILLER_0_129_929 ();
 FILLCELL_X32 FILLER_0_129_961 ();
 FILLCELL_X32 FILLER_0_129_993 ();
 FILLCELL_X32 FILLER_0_129_1025 ();
 FILLCELL_X32 FILLER_0_129_1057 ();
 FILLCELL_X32 FILLER_0_129_1089 ();
 FILLCELL_X16 FILLER_0_129_1121 ();
 FILLCELL_X8 FILLER_0_129_1137 ();
 FILLCELL_X2 FILLER_0_129_1145 ();
 FILLCELL_X1 FILLER_0_129_1147 ();
 FILLCELL_X32 FILLER_0_130_1 ();
 FILLCELL_X32 FILLER_0_130_33 ();
 FILLCELL_X32 FILLER_0_130_65 ();
 FILLCELL_X32 FILLER_0_130_97 ();
 FILLCELL_X32 FILLER_0_130_129 ();
 FILLCELL_X32 FILLER_0_130_161 ();
 FILLCELL_X32 FILLER_0_130_193 ();
 FILLCELL_X32 FILLER_0_130_225 ();
 FILLCELL_X32 FILLER_0_130_257 ();
 FILLCELL_X32 FILLER_0_130_289 ();
 FILLCELL_X32 FILLER_0_130_321 ();
 FILLCELL_X32 FILLER_0_130_353 ();
 FILLCELL_X32 FILLER_0_130_385 ();
 FILLCELL_X32 FILLER_0_130_417 ();
 FILLCELL_X32 FILLER_0_130_449 ();
 FILLCELL_X32 FILLER_0_130_481 ();
 FILLCELL_X32 FILLER_0_130_513 ();
 FILLCELL_X32 FILLER_0_130_545 ();
 FILLCELL_X32 FILLER_0_130_577 ();
 FILLCELL_X16 FILLER_0_130_609 ();
 FILLCELL_X4 FILLER_0_130_625 ();
 FILLCELL_X2 FILLER_0_130_629 ();
 FILLCELL_X32 FILLER_0_130_632 ();
 FILLCELL_X32 FILLER_0_130_664 ();
 FILLCELL_X32 FILLER_0_130_696 ();
 FILLCELL_X32 FILLER_0_130_728 ();
 FILLCELL_X32 FILLER_0_130_760 ();
 FILLCELL_X32 FILLER_0_130_792 ();
 FILLCELL_X32 FILLER_0_130_824 ();
 FILLCELL_X32 FILLER_0_130_856 ();
 FILLCELL_X32 FILLER_0_130_888 ();
 FILLCELL_X32 FILLER_0_130_920 ();
 FILLCELL_X32 FILLER_0_130_952 ();
 FILLCELL_X32 FILLER_0_130_984 ();
 FILLCELL_X32 FILLER_0_130_1016 ();
 FILLCELL_X32 FILLER_0_130_1048 ();
 FILLCELL_X32 FILLER_0_130_1080 ();
 FILLCELL_X32 FILLER_0_130_1112 ();
 FILLCELL_X4 FILLER_0_130_1144 ();
 FILLCELL_X32 FILLER_0_131_1 ();
 FILLCELL_X32 FILLER_0_131_33 ();
 FILLCELL_X32 FILLER_0_131_65 ();
 FILLCELL_X32 FILLER_0_131_97 ();
 FILLCELL_X32 FILLER_0_131_129 ();
 FILLCELL_X32 FILLER_0_131_161 ();
 FILLCELL_X32 FILLER_0_131_193 ();
 FILLCELL_X32 FILLER_0_131_225 ();
 FILLCELL_X32 FILLER_0_131_257 ();
 FILLCELL_X32 FILLER_0_131_289 ();
 FILLCELL_X32 FILLER_0_131_321 ();
 FILLCELL_X32 FILLER_0_131_353 ();
 FILLCELL_X32 FILLER_0_131_385 ();
 FILLCELL_X32 FILLER_0_131_417 ();
 FILLCELL_X32 FILLER_0_131_449 ();
 FILLCELL_X32 FILLER_0_131_481 ();
 FILLCELL_X32 FILLER_0_131_513 ();
 FILLCELL_X32 FILLER_0_131_545 ();
 FILLCELL_X32 FILLER_0_131_577 ();
 FILLCELL_X32 FILLER_0_131_609 ();
 FILLCELL_X32 FILLER_0_131_641 ();
 FILLCELL_X32 FILLER_0_131_673 ();
 FILLCELL_X32 FILLER_0_131_705 ();
 FILLCELL_X32 FILLER_0_131_737 ();
 FILLCELL_X32 FILLER_0_131_769 ();
 FILLCELL_X32 FILLER_0_131_801 ();
 FILLCELL_X32 FILLER_0_131_833 ();
 FILLCELL_X32 FILLER_0_131_865 ();
 FILLCELL_X32 FILLER_0_131_897 ();
 FILLCELL_X32 FILLER_0_131_929 ();
 FILLCELL_X32 FILLER_0_131_961 ();
 FILLCELL_X32 FILLER_0_131_993 ();
 FILLCELL_X32 FILLER_0_131_1025 ();
 FILLCELL_X32 FILLER_0_131_1057 ();
 FILLCELL_X32 FILLER_0_131_1089 ();
 FILLCELL_X16 FILLER_0_131_1121 ();
 FILLCELL_X8 FILLER_0_131_1137 ();
 FILLCELL_X2 FILLER_0_131_1145 ();
 FILLCELL_X1 FILLER_0_131_1147 ();
 FILLCELL_X32 FILLER_0_132_1 ();
 FILLCELL_X32 FILLER_0_132_33 ();
 FILLCELL_X32 FILLER_0_132_65 ();
 FILLCELL_X32 FILLER_0_132_97 ();
 FILLCELL_X32 FILLER_0_132_129 ();
 FILLCELL_X32 FILLER_0_132_161 ();
 FILLCELL_X32 FILLER_0_132_193 ();
 FILLCELL_X32 FILLER_0_132_225 ();
 FILLCELL_X32 FILLER_0_132_257 ();
 FILLCELL_X32 FILLER_0_132_289 ();
 FILLCELL_X32 FILLER_0_132_321 ();
 FILLCELL_X32 FILLER_0_132_353 ();
 FILLCELL_X32 FILLER_0_132_385 ();
 FILLCELL_X32 FILLER_0_132_417 ();
 FILLCELL_X32 FILLER_0_132_449 ();
 FILLCELL_X32 FILLER_0_132_481 ();
 FILLCELL_X32 FILLER_0_132_513 ();
 FILLCELL_X32 FILLER_0_132_545 ();
 FILLCELL_X32 FILLER_0_132_577 ();
 FILLCELL_X16 FILLER_0_132_609 ();
 FILLCELL_X4 FILLER_0_132_625 ();
 FILLCELL_X2 FILLER_0_132_629 ();
 FILLCELL_X32 FILLER_0_132_632 ();
 FILLCELL_X32 FILLER_0_132_664 ();
 FILLCELL_X32 FILLER_0_132_696 ();
 FILLCELL_X32 FILLER_0_132_728 ();
 FILLCELL_X32 FILLER_0_132_760 ();
 FILLCELL_X32 FILLER_0_132_792 ();
 FILLCELL_X32 FILLER_0_132_824 ();
 FILLCELL_X32 FILLER_0_132_856 ();
 FILLCELL_X32 FILLER_0_132_888 ();
 FILLCELL_X32 FILLER_0_132_920 ();
 FILLCELL_X32 FILLER_0_132_952 ();
 FILLCELL_X32 FILLER_0_132_984 ();
 FILLCELL_X32 FILLER_0_132_1016 ();
 FILLCELL_X32 FILLER_0_132_1048 ();
 FILLCELL_X32 FILLER_0_132_1080 ();
 FILLCELL_X32 FILLER_0_132_1112 ();
 FILLCELL_X4 FILLER_0_132_1144 ();
 FILLCELL_X32 FILLER_0_133_1 ();
 FILLCELL_X32 FILLER_0_133_33 ();
 FILLCELL_X32 FILLER_0_133_65 ();
 FILLCELL_X32 FILLER_0_133_97 ();
 FILLCELL_X32 FILLER_0_133_129 ();
 FILLCELL_X32 FILLER_0_133_161 ();
 FILLCELL_X32 FILLER_0_133_193 ();
 FILLCELL_X32 FILLER_0_133_225 ();
 FILLCELL_X32 FILLER_0_133_257 ();
 FILLCELL_X32 FILLER_0_133_289 ();
 FILLCELL_X32 FILLER_0_133_321 ();
 FILLCELL_X32 FILLER_0_133_353 ();
 FILLCELL_X32 FILLER_0_133_385 ();
 FILLCELL_X32 FILLER_0_133_417 ();
 FILLCELL_X32 FILLER_0_133_449 ();
 FILLCELL_X32 FILLER_0_133_481 ();
 FILLCELL_X32 FILLER_0_133_513 ();
 FILLCELL_X32 FILLER_0_133_545 ();
 FILLCELL_X32 FILLER_0_133_577 ();
 FILLCELL_X32 FILLER_0_133_609 ();
 FILLCELL_X32 FILLER_0_133_641 ();
 FILLCELL_X32 FILLER_0_133_673 ();
 FILLCELL_X32 FILLER_0_133_705 ();
 FILLCELL_X32 FILLER_0_133_737 ();
 FILLCELL_X32 FILLER_0_133_769 ();
 FILLCELL_X32 FILLER_0_133_801 ();
 FILLCELL_X32 FILLER_0_133_833 ();
 FILLCELL_X32 FILLER_0_133_865 ();
 FILLCELL_X32 FILLER_0_133_897 ();
 FILLCELL_X32 FILLER_0_133_929 ();
 FILLCELL_X32 FILLER_0_133_961 ();
 FILLCELL_X32 FILLER_0_133_993 ();
 FILLCELL_X32 FILLER_0_133_1025 ();
 FILLCELL_X32 FILLER_0_133_1057 ();
 FILLCELL_X32 FILLER_0_133_1089 ();
 FILLCELL_X16 FILLER_0_133_1121 ();
 FILLCELL_X8 FILLER_0_133_1137 ();
 FILLCELL_X2 FILLER_0_133_1145 ();
 FILLCELL_X1 FILLER_0_133_1147 ();
 FILLCELL_X32 FILLER_0_134_1 ();
 FILLCELL_X32 FILLER_0_134_33 ();
 FILLCELL_X32 FILLER_0_134_65 ();
 FILLCELL_X32 FILLER_0_134_97 ();
 FILLCELL_X32 FILLER_0_134_129 ();
 FILLCELL_X32 FILLER_0_134_161 ();
 FILLCELL_X32 FILLER_0_134_193 ();
 FILLCELL_X32 FILLER_0_134_225 ();
 FILLCELL_X32 FILLER_0_134_257 ();
 FILLCELL_X32 FILLER_0_134_289 ();
 FILLCELL_X32 FILLER_0_134_321 ();
 FILLCELL_X32 FILLER_0_134_353 ();
 FILLCELL_X32 FILLER_0_134_385 ();
 FILLCELL_X32 FILLER_0_134_417 ();
 FILLCELL_X32 FILLER_0_134_449 ();
 FILLCELL_X32 FILLER_0_134_481 ();
 FILLCELL_X32 FILLER_0_134_513 ();
 FILLCELL_X32 FILLER_0_134_545 ();
 FILLCELL_X32 FILLER_0_134_577 ();
 FILLCELL_X16 FILLER_0_134_609 ();
 FILLCELL_X4 FILLER_0_134_625 ();
 FILLCELL_X2 FILLER_0_134_629 ();
 FILLCELL_X32 FILLER_0_134_632 ();
 FILLCELL_X32 FILLER_0_134_664 ();
 FILLCELL_X32 FILLER_0_134_696 ();
 FILLCELL_X32 FILLER_0_134_728 ();
 FILLCELL_X32 FILLER_0_134_760 ();
 FILLCELL_X32 FILLER_0_134_792 ();
 FILLCELL_X32 FILLER_0_134_824 ();
 FILLCELL_X32 FILLER_0_134_856 ();
 FILLCELL_X32 FILLER_0_134_888 ();
 FILLCELL_X32 FILLER_0_134_920 ();
 FILLCELL_X32 FILLER_0_134_952 ();
 FILLCELL_X32 FILLER_0_134_984 ();
 FILLCELL_X32 FILLER_0_134_1016 ();
 FILLCELL_X32 FILLER_0_134_1048 ();
 FILLCELL_X32 FILLER_0_134_1080 ();
 FILLCELL_X32 FILLER_0_134_1112 ();
 FILLCELL_X4 FILLER_0_134_1144 ();
 FILLCELL_X32 FILLER_0_135_1 ();
 FILLCELL_X32 FILLER_0_135_33 ();
 FILLCELL_X32 FILLER_0_135_65 ();
 FILLCELL_X32 FILLER_0_135_97 ();
 FILLCELL_X32 FILLER_0_135_129 ();
 FILLCELL_X32 FILLER_0_135_161 ();
 FILLCELL_X32 FILLER_0_135_193 ();
 FILLCELL_X32 FILLER_0_135_225 ();
 FILLCELL_X32 FILLER_0_135_257 ();
 FILLCELL_X32 FILLER_0_135_289 ();
 FILLCELL_X32 FILLER_0_135_321 ();
 FILLCELL_X32 FILLER_0_135_353 ();
 FILLCELL_X32 FILLER_0_135_385 ();
 FILLCELL_X32 FILLER_0_135_417 ();
 FILLCELL_X32 FILLER_0_135_449 ();
 FILLCELL_X32 FILLER_0_135_481 ();
 FILLCELL_X32 FILLER_0_135_513 ();
 FILLCELL_X32 FILLER_0_135_545 ();
 FILLCELL_X32 FILLER_0_135_577 ();
 FILLCELL_X32 FILLER_0_135_609 ();
 FILLCELL_X32 FILLER_0_135_641 ();
 FILLCELL_X32 FILLER_0_135_673 ();
 FILLCELL_X32 FILLER_0_135_705 ();
 FILLCELL_X32 FILLER_0_135_737 ();
 FILLCELL_X32 FILLER_0_135_769 ();
 FILLCELL_X32 FILLER_0_135_801 ();
 FILLCELL_X32 FILLER_0_135_833 ();
 FILLCELL_X32 FILLER_0_135_865 ();
 FILLCELL_X32 FILLER_0_135_897 ();
 FILLCELL_X32 FILLER_0_135_929 ();
 FILLCELL_X32 FILLER_0_135_961 ();
 FILLCELL_X32 FILLER_0_135_993 ();
 FILLCELL_X32 FILLER_0_135_1025 ();
 FILLCELL_X32 FILLER_0_135_1057 ();
 FILLCELL_X32 FILLER_0_135_1089 ();
 FILLCELL_X16 FILLER_0_135_1121 ();
 FILLCELL_X8 FILLER_0_135_1137 ();
 FILLCELL_X2 FILLER_0_135_1145 ();
 FILLCELL_X1 FILLER_0_135_1147 ();
 FILLCELL_X32 FILLER_0_136_1 ();
 FILLCELL_X32 FILLER_0_136_33 ();
 FILLCELL_X32 FILLER_0_136_65 ();
 FILLCELL_X32 FILLER_0_136_97 ();
 FILLCELL_X32 FILLER_0_136_129 ();
 FILLCELL_X32 FILLER_0_136_161 ();
 FILLCELL_X32 FILLER_0_136_193 ();
 FILLCELL_X32 FILLER_0_136_225 ();
 FILLCELL_X32 FILLER_0_136_257 ();
 FILLCELL_X32 FILLER_0_136_289 ();
 FILLCELL_X32 FILLER_0_136_321 ();
 FILLCELL_X32 FILLER_0_136_353 ();
 FILLCELL_X32 FILLER_0_136_385 ();
 FILLCELL_X32 FILLER_0_136_417 ();
 FILLCELL_X32 FILLER_0_136_449 ();
 FILLCELL_X32 FILLER_0_136_481 ();
 FILLCELL_X32 FILLER_0_136_513 ();
 FILLCELL_X32 FILLER_0_136_545 ();
 FILLCELL_X32 FILLER_0_136_577 ();
 FILLCELL_X16 FILLER_0_136_609 ();
 FILLCELL_X4 FILLER_0_136_625 ();
 FILLCELL_X2 FILLER_0_136_629 ();
 FILLCELL_X32 FILLER_0_136_632 ();
 FILLCELL_X32 FILLER_0_136_664 ();
 FILLCELL_X32 FILLER_0_136_696 ();
 FILLCELL_X32 FILLER_0_136_728 ();
 FILLCELL_X32 FILLER_0_136_760 ();
 FILLCELL_X32 FILLER_0_136_792 ();
 FILLCELL_X32 FILLER_0_136_824 ();
 FILLCELL_X32 FILLER_0_136_856 ();
 FILLCELL_X32 FILLER_0_136_888 ();
 FILLCELL_X32 FILLER_0_136_920 ();
 FILLCELL_X32 FILLER_0_136_952 ();
 FILLCELL_X32 FILLER_0_136_984 ();
 FILLCELL_X32 FILLER_0_136_1016 ();
 FILLCELL_X32 FILLER_0_136_1048 ();
 FILLCELL_X32 FILLER_0_136_1080 ();
 FILLCELL_X32 FILLER_0_136_1112 ();
 FILLCELL_X4 FILLER_0_136_1144 ();
 FILLCELL_X32 FILLER_0_137_1 ();
 FILLCELL_X32 FILLER_0_137_33 ();
 FILLCELL_X32 FILLER_0_137_65 ();
 FILLCELL_X32 FILLER_0_137_97 ();
 FILLCELL_X32 FILLER_0_137_129 ();
 FILLCELL_X32 FILLER_0_137_161 ();
 FILLCELL_X32 FILLER_0_137_193 ();
 FILLCELL_X32 FILLER_0_137_225 ();
 FILLCELL_X32 FILLER_0_137_257 ();
 FILLCELL_X32 FILLER_0_137_289 ();
 FILLCELL_X32 FILLER_0_137_321 ();
 FILLCELL_X32 FILLER_0_137_353 ();
 FILLCELL_X32 FILLER_0_137_385 ();
 FILLCELL_X32 FILLER_0_137_417 ();
 FILLCELL_X32 FILLER_0_137_449 ();
 FILLCELL_X32 FILLER_0_137_481 ();
 FILLCELL_X32 FILLER_0_137_513 ();
 FILLCELL_X32 FILLER_0_137_545 ();
 FILLCELL_X32 FILLER_0_137_577 ();
 FILLCELL_X32 FILLER_0_137_609 ();
 FILLCELL_X32 FILLER_0_137_641 ();
 FILLCELL_X32 FILLER_0_137_673 ();
 FILLCELL_X32 FILLER_0_137_705 ();
 FILLCELL_X32 FILLER_0_137_737 ();
 FILLCELL_X32 FILLER_0_137_769 ();
 FILLCELL_X32 FILLER_0_137_801 ();
 FILLCELL_X32 FILLER_0_137_833 ();
 FILLCELL_X32 FILLER_0_137_865 ();
 FILLCELL_X32 FILLER_0_137_897 ();
 FILLCELL_X32 FILLER_0_137_929 ();
 FILLCELL_X32 FILLER_0_137_961 ();
 FILLCELL_X32 FILLER_0_137_993 ();
 FILLCELL_X32 FILLER_0_137_1025 ();
 FILLCELL_X32 FILLER_0_137_1057 ();
 FILLCELL_X32 FILLER_0_137_1089 ();
 FILLCELL_X16 FILLER_0_137_1121 ();
 FILLCELL_X8 FILLER_0_137_1137 ();
 FILLCELL_X2 FILLER_0_137_1145 ();
 FILLCELL_X1 FILLER_0_137_1147 ();
 FILLCELL_X32 FILLER_0_138_1 ();
 FILLCELL_X32 FILLER_0_138_33 ();
 FILLCELL_X32 FILLER_0_138_65 ();
 FILLCELL_X32 FILLER_0_138_97 ();
 FILLCELL_X32 FILLER_0_138_129 ();
 FILLCELL_X32 FILLER_0_138_161 ();
 FILLCELL_X32 FILLER_0_138_193 ();
 FILLCELL_X32 FILLER_0_138_225 ();
 FILLCELL_X32 FILLER_0_138_257 ();
 FILLCELL_X32 FILLER_0_138_289 ();
 FILLCELL_X32 FILLER_0_138_321 ();
 FILLCELL_X32 FILLER_0_138_353 ();
 FILLCELL_X32 FILLER_0_138_385 ();
 FILLCELL_X32 FILLER_0_138_417 ();
 FILLCELL_X32 FILLER_0_138_449 ();
 FILLCELL_X32 FILLER_0_138_481 ();
 FILLCELL_X32 FILLER_0_138_513 ();
 FILLCELL_X32 FILLER_0_138_545 ();
 FILLCELL_X32 FILLER_0_138_577 ();
 FILLCELL_X16 FILLER_0_138_609 ();
 FILLCELL_X4 FILLER_0_138_625 ();
 FILLCELL_X2 FILLER_0_138_629 ();
 FILLCELL_X32 FILLER_0_138_632 ();
 FILLCELL_X32 FILLER_0_138_664 ();
 FILLCELL_X32 FILLER_0_138_696 ();
 FILLCELL_X32 FILLER_0_138_728 ();
 FILLCELL_X32 FILLER_0_138_760 ();
 FILLCELL_X32 FILLER_0_138_792 ();
 FILLCELL_X32 FILLER_0_138_824 ();
 FILLCELL_X32 FILLER_0_138_856 ();
 FILLCELL_X32 FILLER_0_138_888 ();
 FILLCELL_X32 FILLER_0_138_920 ();
 FILLCELL_X32 FILLER_0_138_952 ();
 FILLCELL_X32 FILLER_0_138_984 ();
 FILLCELL_X32 FILLER_0_138_1016 ();
 FILLCELL_X32 FILLER_0_138_1048 ();
 FILLCELL_X32 FILLER_0_138_1080 ();
 FILLCELL_X32 FILLER_0_138_1112 ();
 FILLCELL_X4 FILLER_0_138_1144 ();
 FILLCELL_X32 FILLER_0_139_1 ();
 FILLCELL_X32 FILLER_0_139_33 ();
 FILLCELL_X32 FILLER_0_139_65 ();
 FILLCELL_X32 FILLER_0_139_97 ();
 FILLCELL_X32 FILLER_0_139_129 ();
 FILLCELL_X32 FILLER_0_139_161 ();
 FILLCELL_X32 FILLER_0_139_193 ();
 FILLCELL_X32 FILLER_0_139_225 ();
 FILLCELL_X32 FILLER_0_139_257 ();
 FILLCELL_X32 FILLER_0_139_289 ();
 FILLCELL_X32 FILLER_0_139_321 ();
 FILLCELL_X32 FILLER_0_139_353 ();
 FILLCELL_X32 FILLER_0_139_385 ();
 FILLCELL_X32 FILLER_0_139_417 ();
 FILLCELL_X32 FILLER_0_139_449 ();
 FILLCELL_X32 FILLER_0_139_481 ();
 FILLCELL_X32 FILLER_0_139_513 ();
 FILLCELL_X32 FILLER_0_139_545 ();
 FILLCELL_X32 FILLER_0_139_577 ();
 FILLCELL_X32 FILLER_0_139_609 ();
 FILLCELL_X32 FILLER_0_139_641 ();
 FILLCELL_X32 FILLER_0_139_673 ();
 FILLCELL_X32 FILLER_0_139_705 ();
 FILLCELL_X32 FILLER_0_139_737 ();
 FILLCELL_X32 FILLER_0_139_769 ();
 FILLCELL_X32 FILLER_0_139_801 ();
 FILLCELL_X32 FILLER_0_139_833 ();
 FILLCELL_X32 FILLER_0_139_865 ();
 FILLCELL_X32 FILLER_0_139_897 ();
 FILLCELL_X32 FILLER_0_139_929 ();
 FILLCELL_X32 FILLER_0_139_961 ();
 FILLCELL_X32 FILLER_0_139_993 ();
 FILLCELL_X32 FILLER_0_139_1025 ();
 FILLCELL_X32 FILLER_0_139_1057 ();
 FILLCELL_X32 FILLER_0_139_1089 ();
 FILLCELL_X16 FILLER_0_139_1121 ();
 FILLCELL_X8 FILLER_0_139_1137 ();
 FILLCELL_X2 FILLER_0_139_1145 ();
 FILLCELL_X1 FILLER_0_139_1147 ();
 FILLCELL_X32 FILLER_0_140_1 ();
 FILLCELL_X32 FILLER_0_140_33 ();
 FILLCELL_X32 FILLER_0_140_65 ();
 FILLCELL_X32 FILLER_0_140_97 ();
 FILLCELL_X32 FILLER_0_140_129 ();
 FILLCELL_X32 FILLER_0_140_161 ();
 FILLCELL_X32 FILLER_0_140_193 ();
 FILLCELL_X32 FILLER_0_140_225 ();
 FILLCELL_X32 FILLER_0_140_257 ();
 FILLCELL_X32 FILLER_0_140_289 ();
 FILLCELL_X32 FILLER_0_140_321 ();
 FILLCELL_X32 FILLER_0_140_353 ();
 FILLCELL_X32 FILLER_0_140_385 ();
 FILLCELL_X32 FILLER_0_140_417 ();
 FILLCELL_X32 FILLER_0_140_449 ();
 FILLCELL_X32 FILLER_0_140_481 ();
 FILLCELL_X32 FILLER_0_140_513 ();
 FILLCELL_X32 FILLER_0_140_545 ();
 FILLCELL_X32 FILLER_0_140_577 ();
 FILLCELL_X16 FILLER_0_140_609 ();
 FILLCELL_X4 FILLER_0_140_625 ();
 FILLCELL_X2 FILLER_0_140_629 ();
 FILLCELL_X32 FILLER_0_140_632 ();
 FILLCELL_X32 FILLER_0_140_664 ();
 FILLCELL_X32 FILLER_0_140_696 ();
 FILLCELL_X32 FILLER_0_140_728 ();
 FILLCELL_X32 FILLER_0_140_760 ();
 FILLCELL_X32 FILLER_0_140_792 ();
 FILLCELL_X32 FILLER_0_140_824 ();
 FILLCELL_X32 FILLER_0_140_856 ();
 FILLCELL_X32 FILLER_0_140_888 ();
 FILLCELL_X32 FILLER_0_140_920 ();
 FILLCELL_X32 FILLER_0_140_952 ();
 FILLCELL_X32 FILLER_0_140_984 ();
 FILLCELL_X32 FILLER_0_140_1016 ();
 FILLCELL_X32 FILLER_0_140_1048 ();
 FILLCELL_X32 FILLER_0_140_1080 ();
 FILLCELL_X32 FILLER_0_140_1112 ();
 FILLCELL_X4 FILLER_0_140_1144 ();
 FILLCELL_X32 FILLER_0_141_1 ();
 FILLCELL_X32 FILLER_0_141_33 ();
 FILLCELL_X32 FILLER_0_141_65 ();
 FILLCELL_X32 FILLER_0_141_97 ();
 FILLCELL_X32 FILLER_0_141_129 ();
 FILLCELL_X32 FILLER_0_141_161 ();
 FILLCELL_X32 FILLER_0_141_193 ();
 FILLCELL_X32 FILLER_0_141_225 ();
 FILLCELL_X32 FILLER_0_141_257 ();
 FILLCELL_X32 FILLER_0_141_289 ();
 FILLCELL_X32 FILLER_0_141_321 ();
 FILLCELL_X32 FILLER_0_141_353 ();
 FILLCELL_X32 FILLER_0_141_385 ();
 FILLCELL_X32 FILLER_0_141_417 ();
 FILLCELL_X32 FILLER_0_141_449 ();
 FILLCELL_X32 FILLER_0_141_481 ();
 FILLCELL_X32 FILLER_0_141_513 ();
 FILLCELL_X32 FILLER_0_141_545 ();
 FILLCELL_X32 FILLER_0_141_577 ();
 FILLCELL_X32 FILLER_0_141_609 ();
 FILLCELL_X32 FILLER_0_141_641 ();
 FILLCELL_X32 FILLER_0_141_673 ();
 FILLCELL_X32 FILLER_0_141_705 ();
 FILLCELL_X32 FILLER_0_141_737 ();
 FILLCELL_X32 FILLER_0_141_769 ();
 FILLCELL_X32 FILLER_0_141_801 ();
 FILLCELL_X32 FILLER_0_141_833 ();
 FILLCELL_X32 FILLER_0_141_865 ();
 FILLCELL_X32 FILLER_0_141_897 ();
 FILLCELL_X32 FILLER_0_141_929 ();
 FILLCELL_X32 FILLER_0_141_961 ();
 FILLCELL_X32 FILLER_0_141_993 ();
 FILLCELL_X32 FILLER_0_141_1025 ();
 FILLCELL_X32 FILLER_0_141_1057 ();
 FILLCELL_X32 FILLER_0_141_1089 ();
 FILLCELL_X16 FILLER_0_141_1121 ();
 FILLCELL_X8 FILLER_0_141_1137 ();
 FILLCELL_X2 FILLER_0_141_1145 ();
 FILLCELL_X1 FILLER_0_141_1147 ();
 FILLCELL_X32 FILLER_0_142_1 ();
 FILLCELL_X32 FILLER_0_142_33 ();
 FILLCELL_X32 FILLER_0_142_65 ();
 FILLCELL_X32 FILLER_0_142_97 ();
 FILLCELL_X32 FILLER_0_142_129 ();
 FILLCELL_X32 FILLER_0_142_161 ();
 FILLCELL_X32 FILLER_0_142_193 ();
 FILLCELL_X32 FILLER_0_142_225 ();
 FILLCELL_X32 FILLER_0_142_257 ();
 FILLCELL_X32 FILLER_0_142_289 ();
 FILLCELL_X32 FILLER_0_142_321 ();
 FILLCELL_X32 FILLER_0_142_353 ();
 FILLCELL_X32 FILLER_0_142_385 ();
 FILLCELL_X32 FILLER_0_142_417 ();
 FILLCELL_X32 FILLER_0_142_449 ();
 FILLCELL_X32 FILLER_0_142_481 ();
 FILLCELL_X32 FILLER_0_142_513 ();
 FILLCELL_X32 FILLER_0_142_545 ();
 FILLCELL_X32 FILLER_0_142_577 ();
 FILLCELL_X16 FILLER_0_142_609 ();
 FILLCELL_X4 FILLER_0_142_625 ();
 FILLCELL_X2 FILLER_0_142_629 ();
 FILLCELL_X32 FILLER_0_142_632 ();
 FILLCELL_X32 FILLER_0_142_664 ();
 FILLCELL_X32 FILLER_0_142_696 ();
 FILLCELL_X32 FILLER_0_142_728 ();
 FILLCELL_X32 FILLER_0_142_760 ();
 FILLCELL_X32 FILLER_0_142_792 ();
 FILLCELL_X32 FILLER_0_142_824 ();
 FILLCELL_X32 FILLER_0_142_856 ();
 FILLCELL_X32 FILLER_0_142_888 ();
 FILLCELL_X32 FILLER_0_142_920 ();
 FILLCELL_X32 FILLER_0_142_952 ();
 FILLCELL_X32 FILLER_0_142_984 ();
 FILLCELL_X32 FILLER_0_142_1016 ();
 FILLCELL_X32 FILLER_0_142_1048 ();
 FILLCELL_X32 FILLER_0_142_1080 ();
 FILLCELL_X32 FILLER_0_142_1112 ();
 FILLCELL_X4 FILLER_0_142_1144 ();
 FILLCELL_X32 FILLER_0_143_1 ();
 FILLCELL_X32 FILLER_0_143_33 ();
 FILLCELL_X32 FILLER_0_143_65 ();
 FILLCELL_X32 FILLER_0_143_97 ();
 FILLCELL_X32 FILLER_0_143_129 ();
 FILLCELL_X32 FILLER_0_143_161 ();
 FILLCELL_X32 FILLER_0_143_193 ();
 FILLCELL_X32 FILLER_0_143_225 ();
 FILLCELL_X32 FILLER_0_143_257 ();
 FILLCELL_X32 FILLER_0_143_289 ();
 FILLCELL_X32 FILLER_0_143_321 ();
 FILLCELL_X32 FILLER_0_143_353 ();
 FILLCELL_X32 FILLER_0_143_385 ();
 FILLCELL_X32 FILLER_0_143_417 ();
 FILLCELL_X32 FILLER_0_143_449 ();
 FILLCELL_X32 FILLER_0_143_481 ();
 FILLCELL_X32 FILLER_0_143_513 ();
 FILLCELL_X32 FILLER_0_143_545 ();
 FILLCELL_X32 FILLER_0_143_577 ();
 FILLCELL_X32 FILLER_0_143_609 ();
 FILLCELL_X32 FILLER_0_143_641 ();
 FILLCELL_X32 FILLER_0_143_673 ();
 FILLCELL_X32 FILLER_0_143_705 ();
 FILLCELL_X32 FILLER_0_143_737 ();
 FILLCELL_X32 FILLER_0_143_769 ();
 FILLCELL_X32 FILLER_0_143_801 ();
 FILLCELL_X32 FILLER_0_143_833 ();
 FILLCELL_X32 FILLER_0_143_865 ();
 FILLCELL_X32 FILLER_0_143_897 ();
 FILLCELL_X32 FILLER_0_143_929 ();
 FILLCELL_X32 FILLER_0_143_961 ();
 FILLCELL_X32 FILLER_0_143_993 ();
 FILLCELL_X32 FILLER_0_143_1025 ();
 FILLCELL_X32 FILLER_0_143_1057 ();
 FILLCELL_X32 FILLER_0_143_1089 ();
 FILLCELL_X16 FILLER_0_143_1121 ();
 FILLCELL_X8 FILLER_0_143_1137 ();
 FILLCELL_X2 FILLER_0_143_1145 ();
 FILLCELL_X1 FILLER_0_143_1147 ();
 FILLCELL_X32 FILLER_0_144_1 ();
 FILLCELL_X32 FILLER_0_144_33 ();
 FILLCELL_X32 FILLER_0_144_65 ();
 FILLCELL_X32 FILLER_0_144_97 ();
 FILLCELL_X32 FILLER_0_144_129 ();
 FILLCELL_X32 FILLER_0_144_161 ();
 FILLCELL_X32 FILLER_0_144_193 ();
 FILLCELL_X32 FILLER_0_144_225 ();
 FILLCELL_X32 FILLER_0_144_257 ();
 FILLCELL_X32 FILLER_0_144_289 ();
 FILLCELL_X32 FILLER_0_144_321 ();
 FILLCELL_X32 FILLER_0_144_353 ();
 FILLCELL_X32 FILLER_0_144_385 ();
 FILLCELL_X32 FILLER_0_144_417 ();
 FILLCELL_X32 FILLER_0_144_449 ();
 FILLCELL_X32 FILLER_0_144_481 ();
 FILLCELL_X32 FILLER_0_144_513 ();
 FILLCELL_X32 FILLER_0_144_545 ();
 FILLCELL_X32 FILLER_0_144_577 ();
 FILLCELL_X16 FILLER_0_144_609 ();
 FILLCELL_X4 FILLER_0_144_625 ();
 FILLCELL_X2 FILLER_0_144_629 ();
 FILLCELL_X32 FILLER_0_144_632 ();
 FILLCELL_X32 FILLER_0_144_664 ();
 FILLCELL_X32 FILLER_0_144_696 ();
 FILLCELL_X32 FILLER_0_144_728 ();
 FILLCELL_X32 FILLER_0_144_760 ();
 FILLCELL_X32 FILLER_0_144_792 ();
 FILLCELL_X32 FILLER_0_144_824 ();
 FILLCELL_X32 FILLER_0_144_856 ();
 FILLCELL_X32 FILLER_0_144_888 ();
 FILLCELL_X32 FILLER_0_144_920 ();
 FILLCELL_X32 FILLER_0_144_952 ();
 FILLCELL_X32 FILLER_0_144_984 ();
 FILLCELL_X32 FILLER_0_144_1016 ();
 FILLCELL_X32 FILLER_0_144_1048 ();
 FILLCELL_X32 FILLER_0_144_1080 ();
 FILLCELL_X32 FILLER_0_144_1112 ();
 FILLCELL_X4 FILLER_0_144_1144 ();
 FILLCELL_X32 FILLER_0_145_1 ();
 FILLCELL_X32 FILLER_0_145_33 ();
 FILLCELL_X32 FILLER_0_145_65 ();
 FILLCELL_X32 FILLER_0_145_97 ();
 FILLCELL_X32 FILLER_0_145_129 ();
 FILLCELL_X32 FILLER_0_145_161 ();
 FILLCELL_X32 FILLER_0_145_193 ();
 FILLCELL_X32 FILLER_0_145_225 ();
 FILLCELL_X32 FILLER_0_145_257 ();
 FILLCELL_X32 FILLER_0_145_289 ();
 FILLCELL_X32 FILLER_0_145_321 ();
 FILLCELL_X32 FILLER_0_145_353 ();
 FILLCELL_X32 FILLER_0_145_385 ();
 FILLCELL_X32 FILLER_0_145_417 ();
 FILLCELL_X32 FILLER_0_145_449 ();
 FILLCELL_X32 FILLER_0_145_481 ();
 FILLCELL_X32 FILLER_0_145_513 ();
 FILLCELL_X32 FILLER_0_145_545 ();
 FILLCELL_X32 FILLER_0_145_577 ();
 FILLCELL_X32 FILLER_0_145_609 ();
 FILLCELL_X32 FILLER_0_145_641 ();
 FILLCELL_X32 FILLER_0_145_673 ();
 FILLCELL_X32 FILLER_0_145_705 ();
 FILLCELL_X32 FILLER_0_145_737 ();
 FILLCELL_X32 FILLER_0_145_769 ();
 FILLCELL_X32 FILLER_0_145_801 ();
 FILLCELL_X32 FILLER_0_145_833 ();
 FILLCELL_X32 FILLER_0_145_865 ();
 FILLCELL_X32 FILLER_0_145_897 ();
 FILLCELL_X32 FILLER_0_145_929 ();
 FILLCELL_X32 FILLER_0_145_961 ();
 FILLCELL_X32 FILLER_0_145_993 ();
 FILLCELL_X32 FILLER_0_145_1025 ();
 FILLCELL_X32 FILLER_0_145_1057 ();
 FILLCELL_X32 FILLER_0_145_1089 ();
 FILLCELL_X16 FILLER_0_145_1121 ();
 FILLCELL_X8 FILLER_0_145_1137 ();
 FILLCELL_X2 FILLER_0_145_1145 ();
 FILLCELL_X1 FILLER_0_145_1147 ();
 FILLCELL_X32 FILLER_0_146_1 ();
 FILLCELL_X32 FILLER_0_146_33 ();
 FILLCELL_X32 FILLER_0_146_65 ();
 FILLCELL_X32 FILLER_0_146_97 ();
 FILLCELL_X32 FILLER_0_146_129 ();
 FILLCELL_X32 FILLER_0_146_161 ();
 FILLCELL_X32 FILLER_0_146_193 ();
 FILLCELL_X32 FILLER_0_146_225 ();
 FILLCELL_X32 FILLER_0_146_257 ();
 FILLCELL_X32 FILLER_0_146_289 ();
 FILLCELL_X32 FILLER_0_146_321 ();
 FILLCELL_X32 FILLER_0_146_353 ();
 FILLCELL_X32 FILLER_0_146_385 ();
 FILLCELL_X32 FILLER_0_146_417 ();
 FILLCELL_X32 FILLER_0_146_449 ();
 FILLCELL_X32 FILLER_0_146_481 ();
 FILLCELL_X32 FILLER_0_146_513 ();
 FILLCELL_X32 FILLER_0_146_545 ();
 FILLCELL_X32 FILLER_0_146_577 ();
 FILLCELL_X16 FILLER_0_146_609 ();
 FILLCELL_X4 FILLER_0_146_625 ();
 FILLCELL_X2 FILLER_0_146_629 ();
 FILLCELL_X32 FILLER_0_146_632 ();
 FILLCELL_X32 FILLER_0_146_664 ();
 FILLCELL_X32 FILLER_0_146_696 ();
 FILLCELL_X32 FILLER_0_146_728 ();
 FILLCELL_X32 FILLER_0_146_760 ();
 FILLCELL_X32 FILLER_0_146_792 ();
 FILLCELL_X32 FILLER_0_146_824 ();
 FILLCELL_X32 FILLER_0_146_856 ();
 FILLCELL_X32 FILLER_0_146_888 ();
 FILLCELL_X32 FILLER_0_146_920 ();
 FILLCELL_X32 FILLER_0_146_952 ();
 FILLCELL_X32 FILLER_0_146_984 ();
 FILLCELL_X32 FILLER_0_146_1016 ();
 FILLCELL_X32 FILLER_0_146_1048 ();
 FILLCELL_X32 FILLER_0_146_1080 ();
 FILLCELL_X32 FILLER_0_146_1112 ();
 FILLCELL_X4 FILLER_0_146_1144 ();
 FILLCELL_X32 FILLER_0_147_1 ();
 FILLCELL_X32 FILLER_0_147_33 ();
 FILLCELL_X32 FILLER_0_147_65 ();
 FILLCELL_X32 FILLER_0_147_97 ();
 FILLCELL_X32 FILLER_0_147_129 ();
 FILLCELL_X32 FILLER_0_147_161 ();
 FILLCELL_X32 FILLER_0_147_193 ();
 FILLCELL_X32 FILLER_0_147_225 ();
 FILLCELL_X32 FILLER_0_147_257 ();
 FILLCELL_X32 FILLER_0_147_289 ();
 FILLCELL_X32 FILLER_0_147_321 ();
 FILLCELL_X32 FILLER_0_147_353 ();
 FILLCELL_X32 FILLER_0_147_385 ();
 FILLCELL_X32 FILLER_0_147_417 ();
 FILLCELL_X32 FILLER_0_147_449 ();
 FILLCELL_X32 FILLER_0_147_481 ();
 FILLCELL_X32 FILLER_0_147_513 ();
 FILLCELL_X32 FILLER_0_147_545 ();
 FILLCELL_X32 FILLER_0_147_577 ();
 FILLCELL_X32 FILLER_0_147_609 ();
 FILLCELL_X32 FILLER_0_147_641 ();
 FILLCELL_X32 FILLER_0_147_673 ();
 FILLCELL_X32 FILLER_0_147_705 ();
 FILLCELL_X32 FILLER_0_147_737 ();
 FILLCELL_X32 FILLER_0_147_769 ();
 FILLCELL_X32 FILLER_0_147_801 ();
 FILLCELL_X32 FILLER_0_147_833 ();
 FILLCELL_X32 FILLER_0_147_865 ();
 FILLCELL_X32 FILLER_0_147_897 ();
 FILLCELL_X32 FILLER_0_147_929 ();
 FILLCELL_X32 FILLER_0_147_961 ();
 FILLCELL_X32 FILLER_0_147_993 ();
 FILLCELL_X32 FILLER_0_147_1025 ();
 FILLCELL_X32 FILLER_0_147_1057 ();
 FILLCELL_X32 FILLER_0_147_1089 ();
 FILLCELL_X16 FILLER_0_147_1121 ();
 FILLCELL_X8 FILLER_0_147_1137 ();
 FILLCELL_X2 FILLER_0_147_1145 ();
 FILLCELL_X1 FILLER_0_147_1147 ();
 FILLCELL_X32 FILLER_0_148_1 ();
 FILLCELL_X32 FILLER_0_148_33 ();
 FILLCELL_X32 FILLER_0_148_65 ();
 FILLCELL_X32 FILLER_0_148_97 ();
 FILLCELL_X32 FILLER_0_148_129 ();
 FILLCELL_X32 FILLER_0_148_161 ();
 FILLCELL_X32 FILLER_0_148_193 ();
 FILLCELL_X32 FILLER_0_148_225 ();
 FILLCELL_X32 FILLER_0_148_257 ();
 FILLCELL_X32 FILLER_0_148_289 ();
 FILLCELL_X32 FILLER_0_148_321 ();
 FILLCELL_X32 FILLER_0_148_353 ();
 FILLCELL_X32 FILLER_0_148_385 ();
 FILLCELL_X32 FILLER_0_148_417 ();
 FILLCELL_X32 FILLER_0_148_449 ();
 FILLCELL_X32 FILLER_0_148_481 ();
 FILLCELL_X32 FILLER_0_148_513 ();
 FILLCELL_X32 FILLER_0_148_545 ();
 FILLCELL_X32 FILLER_0_148_577 ();
 FILLCELL_X16 FILLER_0_148_609 ();
 FILLCELL_X4 FILLER_0_148_625 ();
 FILLCELL_X2 FILLER_0_148_629 ();
 FILLCELL_X32 FILLER_0_148_632 ();
 FILLCELL_X32 FILLER_0_148_664 ();
 FILLCELL_X32 FILLER_0_148_696 ();
 FILLCELL_X32 FILLER_0_148_728 ();
 FILLCELL_X32 FILLER_0_148_760 ();
 FILLCELL_X32 FILLER_0_148_792 ();
 FILLCELL_X32 FILLER_0_148_824 ();
 FILLCELL_X32 FILLER_0_148_856 ();
 FILLCELL_X32 FILLER_0_148_888 ();
 FILLCELL_X32 FILLER_0_148_920 ();
 FILLCELL_X32 FILLER_0_148_952 ();
 FILLCELL_X32 FILLER_0_148_984 ();
 FILLCELL_X32 FILLER_0_148_1016 ();
 FILLCELL_X32 FILLER_0_148_1048 ();
 FILLCELL_X32 FILLER_0_148_1080 ();
 FILLCELL_X32 FILLER_0_148_1112 ();
 FILLCELL_X4 FILLER_0_148_1144 ();
 FILLCELL_X32 FILLER_0_149_1 ();
 FILLCELL_X32 FILLER_0_149_33 ();
 FILLCELL_X32 FILLER_0_149_65 ();
 FILLCELL_X32 FILLER_0_149_97 ();
 FILLCELL_X32 FILLER_0_149_129 ();
 FILLCELL_X32 FILLER_0_149_161 ();
 FILLCELL_X32 FILLER_0_149_193 ();
 FILLCELL_X32 FILLER_0_149_225 ();
 FILLCELL_X32 FILLER_0_149_257 ();
 FILLCELL_X32 FILLER_0_149_289 ();
 FILLCELL_X32 FILLER_0_149_321 ();
 FILLCELL_X32 FILLER_0_149_353 ();
 FILLCELL_X32 FILLER_0_149_385 ();
 FILLCELL_X32 FILLER_0_149_417 ();
 FILLCELL_X32 FILLER_0_149_449 ();
 FILLCELL_X32 FILLER_0_149_481 ();
 FILLCELL_X32 FILLER_0_149_513 ();
 FILLCELL_X32 FILLER_0_149_545 ();
 FILLCELL_X32 FILLER_0_149_577 ();
 FILLCELL_X32 FILLER_0_149_609 ();
 FILLCELL_X32 FILLER_0_149_641 ();
 FILLCELL_X32 FILLER_0_149_673 ();
 FILLCELL_X32 FILLER_0_149_705 ();
 FILLCELL_X32 FILLER_0_149_737 ();
 FILLCELL_X32 FILLER_0_149_769 ();
 FILLCELL_X32 FILLER_0_149_801 ();
 FILLCELL_X32 FILLER_0_149_833 ();
 FILLCELL_X32 FILLER_0_149_865 ();
 FILLCELL_X32 FILLER_0_149_897 ();
 FILLCELL_X32 FILLER_0_149_929 ();
 FILLCELL_X32 FILLER_0_149_961 ();
 FILLCELL_X32 FILLER_0_149_993 ();
 FILLCELL_X32 FILLER_0_149_1025 ();
 FILLCELL_X32 FILLER_0_149_1057 ();
 FILLCELL_X32 FILLER_0_149_1089 ();
 FILLCELL_X16 FILLER_0_149_1121 ();
 FILLCELL_X8 FILLER_0_149_1137 ();
 FILLCELL_X2 FILLER_0_149_1145 ();
 FILLCELL_X1 FILLER_0_149_1147 ();
 FILLCELL_X32 FILLER_0_150_1 ();
 FILLCELL_X32 FILLER_0_150_33 ();
 FILLCELL_X32 FILLER_0_150_65 ();
 FILLCELL_X32 FILLER_0_150_97 ();
 FILLCELL_X32 FILLER_0_150_129 ();
 FILLCELL_X32 FILLER_0_150_161 ();
 FILLCELL_X32 FILLER_0_150_193 ();
 FILLCELL_X32 FILLER_0_150_225 ();
 FILLCELL_X32 FILLER_0_150_257 ();
 FILLCELL_X32 FILLER_0_150_289 ();
 FILLCELL_X32 FILLER_0_150_321 ();
 FILLCELL_X32 FILLER_0_150_353 ();
 FILLCELL_X32 FILLER_0_150_385 ();
 FILLCELL_X32 FILLER_0_150_417 ();
 FILLCELL_X32 FILLER_0_150_449 ();
 FILLCELL_X32 FILLER_0_150_481 ();
 FILLCELL_X32 FILLER_0_150_513 ();
 FILLCELL_X32 FILLER_0_150_545 ();
 FILLCELL_X32 FILLER_0_150_577 ();
 FILLCELL_X16 FILLER_0_150_609 ();
 FILLCELL_X4 FILLER_0_150_625 ();
 FILLCELL_X2 FILLER_0_150_629 ();
 FILLCELL_X32 FILLER_0_150_632 ();
 FILLCELL_X32 FILLER_0_150_664 ();
 FILLCELL_X32 FILLER_0_150_696 ();
 FILLCELL_X32 FILLER_0_150_728 ();
 FILLCELL_X32 FILLER_0_150_760 ();
 FILLCELL_X32 FILLER_0_150_792 ();
 FILLCELL_X32 FILLER_0_150_824 ();
 FILLCELL_X32 FILLER_0_150_856 ();
 FILLCELL_X32 FILLER_0_150_888 ();
 FILLCELL_X32 FILLER_0_150_920 ();
 FILLCELL_X32 FILLER_0_150_952 ();
 FILLCELL_X32 FILLER_0_150_984 ();
 FILLCELL_X32 FILLER_0_150_1016 ();
 FILLCELL_X32 FILLER_0_150_1048 ();
 FILLCELL_X32 FILLER_0_150_1080 ();
 FILLCELL_X32 FILLER_0_150_1112 ();
 FILLCELL_X4 FILLER_0_150_1144 ();
 FILLCELL_X32 FILLER_0_151_1 ();
 FILLCELL_X32 FILLER_0_151_33 ();
 FILLCELL_X32 FILLER_0_151_65 ();
 FILLCELL_X32 FILLER_0_151_97 ();
 FILLCELL_X32 FILLER_0_151_129 ();
 FILLCELL_X32 FILLER_0_151_161 ();
 FILLCELL_X32 FILLER_0_151_193 ();
 FILLCELL_X32 FILLER_0_151_225 ();
 FILLCELL_X32 FILLER_0_151_257 ();
 FILLCELL_X32 FILLER_0_151_289 ();
 FILLCELL_X32 FILLER_0_151_321 ();
 FILLCELL_X32 FILLER_0_151_353 ();
 FILLCELL_X32 FILLER_0_151_385 ();
 FILLCELL_X32 FILLER_0_151_417 ();
 FILLCELL_X32 FILLER_0_151_449 ();
 FILLCELL_X32 FILLER_0_151_481 ();
 FILLCELL_X32 FILLER_0_151_513 ();
 FILLCELL_X32 FILLER_0_151_545 ();
 FILLCELL_X32 FILLER_0_151_577 ();
 FILLCELL_X32 FILLER_0_151_609 ();
 FILLCELL_X32 FILLER_0_151_641 ();
 FILLCELL_X32 FILLER_0_151_673 ();
 FILLCELL_X32 FILLER_0_151_705 ();
 FILLCELL_X32 FILLER_0_151_737 ();
 FILLCELL_X32 FILLER_0_151_769 ();
 FILLCELL_X32 FILLER_0_151_801 ();
 FILLCELL_X32 FILLER_0_151_833 ();
 FILLCELL_X32 FILLER_0_151_865 ();
 FILLCELL_X32 FILLER_0_151_897 ();
 FILLCELL_X32 FILLER_0_151_929 ();
 FILLCELL_X32 FILLER_0_151_961 ();
 FILLCELL_X32 FILLER_0_151_993 ();
 FILLCELL_X32 FILLER_0_151_1025 ();
 FILLCELL_X32 FILLER_0_151_1057 ();
 FILLCELL_X32 FILLER_0_151_1089 ();
 FILLCELL_X16 FILLER_0_151_1121 ();
 FILLCELL_X8 FILLER_0_151_1137 ();
 FILLCELL_X2 FILLER_0_151_1145 ();
 FILLCELL_X1 FILLER_0_151_1147 ();
 FILLCELL_X32 FILLER_0_152_1 ();
 FILLCELL_X32 FILLER_0_152_33 ();
 FILLCELL_X32 FILLER_0_152_65 ();
 FILLCELL_X32 FILLER_0_152_97 ();
 FILLCELL_X32 FILLER_0_152_129 ();
 FILLCELL_X32 FILLER_0_152_161 ();
 FILLCELL_X32 FILLER_0_152_193 ();
 FILLCELL_X32 FILLER_0_152_225 ();
 FILLCELL_X32 FILLER_0_152_257 ();
 FILLCELL_X32 FILLER_0_152_289 ();
 FILLCELL_X32 FILLER_0_152_321 ();
 FILLCELL_X32 FILLER_0_152_353 ();
 FILLCELL_X32 FILLER_0_152_385 ();
 FILLCELL_X32 FILLER_0_152_417 ();
 FILLCELL_X32 FILLER_0_152_449 ();
 FILLCELL_X32 FILLER_0_152_481 ();
 FILLCELL_X32 FILLER_0_152_513 ();
 FILLCELL_X32 FILLER_0_152_545 ();
 FILLCELL_X32 FILLER_0_152_577 ();
 FILLCELL_X16 FILLER_0_152_609 ();
 FILLCELL_X4 FILLER_0_152_625 ();
 FILLCELL_X2 FILLER_0_152_629 ();
 FILLCELL_X32 FILLER_0_152_632 ();
 FILLCELL_X32 FILLER_0_152_664 ();
 FILLCELL_X32 FILLER_0_152_696 ();
 FILLCELL_X32 FILLER_0_152_728 ();
 FILLCELL_X32 FILLER_0_152_760 ();
 FILLCELL_X32 FILLER_0_152_792 ();
 FILLCELL_X32 FILLER_0_152_824 ();
 FILLCELL_X32 FILLER_0_152_856 ();
 FILLCELL_X32 FILLER_0_152_888 ();
 FILLCELL_X32 FILLER_0_152_920 ();
 FILLCELL_X32 FILLER_0_152_952 ();
 FILLCELL_X32 FILLER_0_152_984 ();
 FILLCELL_X32 FILLER_0_152_1016 ();
 FILLCELL_X32 FILLER_0_152_1048 ();
 FILLCELL_X32 FILLER_0_152_1080 ();
 FILLCELL_X32 FILLER_0_152_1112 ();
 FILLCELL_X4 FILLER_0_152_1144 ();
 FILLCELL_X32 FILLER_0_153_1 ();
 FILLCELL_X32 FILLER_0_153_33 ();
 FILLCELL_X32 FILLER_0_153_65 ();
 FILLCELL_X32 FILLER_0_153_97 ();
 FILLCELL_X32 FILLER_0_153_129 ();
 FILLCELL_X32 FILLER_0_153_161 ();
 FILLCELL_X32 FILLER_0_153_193 ();
 FILLCELL_X32 FILLER_0_153_225 ();
 FILLCELL_X32 FILLER_0_153_257 ();
 FILLCELL_X32 FILLER_0_153_289 ();
 FILLCELL_X32 FILLER_0_153_321 ();
 FILLCELL_X32 FILLER_0_153_353 ();
 FILLCELL_X32 FILLER_0_153_385 ();
 FILLCELL_X32 FILLER_0_153_417 ();
 FILLCELL_X32 FILLER_0_153_449 ();
 FILLCELL_X32 FILLER_0_153_481 ();
 FILLCELL_X32 FILLER_0_153_513 ();
 FILLCELL_X32 FILLER_0_153_545 ();
 FILLCELL_X32 FILLER_0_153_577 ();
 FILLCELL_X32 FILLER_0_153_609 ();
 FILLCELL_X32 FILLER_0_153_641 ();
 FILLCELL_X32 FILLER_0_153_673 ();
 FILLCELL_X32 FILLER_0_153_705 ();
 FILLCELL_X32 FILLER_0_153_737 ();
 FILLCELL_X32 FILLER_0_153_769 ();
 FILLCELL_X32 FILLER_0_153_801 ();
 FILLCELL_X32 FILLER_0_153_833 ();
 FILLCELL_X32 FILLER_0_153_865 ();
 FILLCELL_X32 FILLER_0_153_897 ();
 FILLCELL_X32 FILLER_0_153_929 ();
 FILLCELL_X32 FILLER_0_153_961 ();
 FILLCELL_X32 FILLER_0_153_993 ();
 FILLCELL_X32 FILLER_0_153_1025 ();
 FILLCELL_X32 FILLER_0_153_1057 ();
 FILLCELL_X32 FILLER_0_153_1089 ();
 FILLCELL_X16 FILLER_0_153_1121 ();
 FILLCELL_X8 FILLER_0_153_1137 ();
 FILLCELL_X2 FILLER_0_153_1145 ();
 FILLCELL_X1 FILLER_0_153_1147 ();
 FILLCELL_X32 FILLER_0_154_1 ();
 FILLCELL_X32 FILLER_0_154_33 ();
 FILLCELL_X32 FILLER_0_154_65 ();
 FILLCELL_X32 FILLER_0_154_97 ();
 FILLCELL_X32 FILLER_0_154_129 ();
 FILLCELL_X32 FILLER_0_154_161 ();
 FILLCELL_X32 FILLER_0_154_193 ();
 FILLCELL_X32 FILLER_0_154_225 ();
 FILLCELL_X32 FILLER_0_154_257 ();
 FILLCELL_X32 FILLER_0_154_289 ();
 FILLCELL_X32 FILLER_0_154_321 ();
 FILLCELL_X32 FILLER_0_154_353 ();
 FILLCELL_X32 FILLER_0_154_385 ();
 FILLCELL_X32 FILLER_0_154_417 ();
 FILLCELL_X32 FILLER_0_154_449 ();
 FILLCELL_X32 FILLER_0_154_481 ();
 FILLCELL_X32 FILLER_0_154_513 ();
 FILLCELL_X32 FILLER_0_154_545 ();
 FILLCELL_X32 FILLER_0_154_577 ();
 FILLCELL_X16 FILLER_0_154_609 ();
 FILLCELL_X4 FILLER_0_154_625 ();
 FILLCELL_X2 FILLER_0_154_629 ();
 FILLCELL_X32 FILLER_0_154_632 ();
 FILLCELL_X32 FILLER_0_154_664 ();
 FILLCELL_X32 FILLER_0_154_696 ();
 FILLCELL_X32 FILLER_0_154_728 ();
 FILLCELL_X32 FILLER_0_154_760 ();
 FILLCELL_X32 FILLER_0_154_792 ();
 FILLCELL_X32 FILLER_0_154_824 ();
 FILLCELL_X32 FILLER_0_154_856 ();
 FILLCELL_X32 FILLER_0_154_888 ();
 FILLCELL_X32 FILLER_0_154_920 ();
 FILLCELL_X32 FILLER_0_154_952 ();
 FILLCELL_X32 FILLER_0_154_984 ();
 FILLCELL_X32 FILLER_0_154_1016 ();
 FILLCELL_X32 FILLER_0_154_1048 ();
 FILLCELL_X32 FILLER_0_154_1080 ();
 FILLCELL_X32 FILLER_0_154_1112 ();
 FILLCELL_X4 FILLER_0_154_1144 ();
endmodule
